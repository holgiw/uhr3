PK
     ���Z�ަ���  ��     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_0":[],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_1":["pin-type-component_b21448dd-3ab4-402c-a381-8ae77300b5cc_1"],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_2":["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_0"],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_3":["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_4"],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_4":[],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_5":["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_3"],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_6":["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_1"],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_7":["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_6","pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_1"],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_8":["pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_0"],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_9":["pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_1"],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_10":["pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_1"],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_11":[],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_12":[],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_13":[],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_14":[],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_15":[],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_16":[],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_17":["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_5"],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_18":["pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_2"],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_19":[],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_20":["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_2"],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_21":[],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_22":[],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_23":[],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_24":[],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_25":[],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_26":[],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_27":[],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_28":[],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_29":[],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_30":[],"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_31":[],"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_0":["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_2"],"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_1":["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_6"],"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_2":["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_20"],"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_3":["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_5"],"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_4":["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_3"],"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_5":["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_17"],"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_6":["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_7"],"pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_0":["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_8"],"pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_1":["pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_0","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_9"],"pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_0":["pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_1","pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_0"],"pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_1":["pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_1","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_10"],"pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_0":["pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_0"],"pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_1":["pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_1"],"pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_0":[],"pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_1":["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_7"],"pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_2":["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_18"],"pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_3":[],"pin-type-component_b21448dd-3ab4-402c-a381-8ae77300b5cc_0":[],"pin-type-component_b21448dd-3ab4-402c-a381-8ae77300b5cc_1":["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_1"]},"pin_to_color":{"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_0":"#000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_1":"#C28C9F","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_2":"#804040","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_3":"#FFE502","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_4":"#000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_5":"#005F39","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_6":"#ffffff","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_7":"#ff0000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_8":"#c0c0c0","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_9":"#c0c0c0","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_10":"#c0c0c0","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_11":"#000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_12":"#000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_13":"#000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_14":"#000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_15":"#000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_16":"#000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_17":"#0080ff","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_18":"#00AE7E","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_19":"#000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_20":"#ff8000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_21":"#000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_22":"#000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_23":"#000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_24":"#000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_25":"#000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_26":"#000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_27":"#000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_28":"#000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_29":"#000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_30":"#000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_31":"#000000","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_0":"#804040","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_1":"#ffffff","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_2":"#ff8000","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_3":"#005F39","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_4":"#FFE502","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_5":"#0080ff","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_6":"#ff0000","pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_0":"#c0c0c0","pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_1":"#c0c0c0","pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_0":"#c0c0c0","pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_1":"#c0c0c0","pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_0":"#c0c0c0","pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_1":"#c0c0c0","pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_0":"#000000","pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_1":"#ff0000","pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_2":"#00AE7E","pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_3":"#000000","pin-type-component_b21448dd-3ab4-402c-a381-8ae77300b5cc_0":"#000000","pin-type-component_b21448dd-3ab4-402c-a381-8ae77300b5cc_1":"#C28C9F"},"pin_to_state":{"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_0":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_1":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_2":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_3":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_4":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_5":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_6":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_7":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_8":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_9":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_10":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_11":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_12":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_13":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_14":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_15":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_16":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_17":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_18":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_19":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_20":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_21":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_22":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_23":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_24":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_25":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_26":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_27":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_28":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_29":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_30":"neutral","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_31":"neutral","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_0":"neutral","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_1":"neutral","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_2":"neutral","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_3":"neutral","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_4":"neutral","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_5":"neutral","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_6":"neutral","pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_0":"neutral","pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_1":"neutral","pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_0":"neutral","pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_1":"neutral","pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_0":"neutral","pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_1":"neutral","pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_0":"neutral","pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_1":"neutral","pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_2":"neutral","pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_3":"neutral","pin-type-component_b21448dd-3ab4-402c-a381-8ae77300b5cc_0":"neutral","pin-type-component_b21448dd-3ab4-402c-a381-8ae77300b5cc_1":"neutral"},"next_color_idx":13,"wires_placed_in_order":[["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_7","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_6"],["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_17","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_5"],["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_2","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_20"],["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_4","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_3"],["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_3","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_5"],["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_1","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_6"],["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_0","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_2"],["pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_0","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_23"],["pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_1","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_22"],["pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_1","pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_0"],["pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_1","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_21"],["pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_0","pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_0"],["pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_1","pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_1"],["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_8","pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_0"],["pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_1","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_9"],["pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_1","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_10"],["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_18","pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_2"],["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_7","pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_1"],["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_1","pin-type-component_b21448dd-3ab4-402c-a381-8ae77300b5cc_1"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_7","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_6"]]],[[],[["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_17","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_5"]]],[[],[["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_2","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_20"]]],[[],[["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_4","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_3"]]],[[],[["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_3","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_5"]]],[[],[["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_1","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_6"]]],[[],[["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_0","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_2"]]],[[],[["pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_0","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_23"]]],[[],[["pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_1","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_22"]]],[[],[["pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_1","pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_0"]]],[[],[["pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_1","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_21"]]],[[],[["pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_0","pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_0"]]],[[],[["pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_1","pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_1"]]],[[["pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_0","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_23"]],[]],[[["pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_1","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_22"]],[]],[[["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_21","pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_1"]],[]],[[],[["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_8","pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_0"]]],[[],[["pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_1","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_9"]]],[[],[["pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_1","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_10"]]],[[],[["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_18","pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_2"]]],[[],[["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_7","pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_1"]]],[[],[["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_1","pin-type-component_b21448dd-3ab4-402c-a381-8ae77300b5cc_1"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_0":"_","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_1":"0000000000000011","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_2":"0000000000000006","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_3":"0000000000000003","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_4":"_","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_5":"0000000000000004","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_6":"0000000000000005","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_7":"0000000000000000","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_8":"0000000000000007","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_9":"0000000000000008","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_10":"0000000000000009","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_11":"_","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_12":"_","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_13":"_","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_14":"_","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_15":"_","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_16":"_","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_17":"0000000000000001","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_18":"0000000000000010","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_19":"_","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_20":"0000000000000002","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_21":"_","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_22":"_","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_23":"_","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_24":"_","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_25":"_","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_26":"_","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_27":"_","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_28":"_","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_29":"_","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_30":"_","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_31":"_","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_0":"0000000000000006","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_1":"0000000000000005","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_2":"0000000000000002","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_3":"0000000000000004","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_4":"0000000000000003","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_5":"0000000000000001","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_6":"0000000000000000","pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_0":"0000000000000007","pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_1":"0000000000000008","pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_0":"0000000000000008","pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_1":"0000000000000009","pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_0":"0000000000000008","pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_1":"0000000000000009","pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_0":"_","pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_1":"0000000000000000","pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_2":"0000000000000010","pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_3":"_","pin-type-component_b21448dd-3ab4-402c-a381-8ae77300b5cc_0":"_","pin-type-component_b21448dd-3ab4-402c-a381-8ae77300b5cc_1":"0000000000000011"},"component_id_to_pins":{"aff8a528-b934-4625-84af-01f958e4a790":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31"],"41fc28b8-a12b-46bf-af23-3da2617c8a06":["0","1","2","3","4","5","6"],"20642084-3e38-42a8-864e-12f237eae7bb":["0","1"],"e95d33f2-d715-46ec-8052-7ee80f0ef8db":["0","1"],"07565f67-0738-4731-9f74-672de39f4e2e":["0","1"],"c658a115-ed11-4c13-aea5-34348036d108":["0","1","2","3"],"96dc7d5d-837f-47c8-b317-a9d24f1c8303":[],"89c3afb5-35ce-4fba-a71b-117023af28ae":[],"ede89323-f462-4ac4-a580-8d3a6368b911":[],"b21448dd-3ab4-402c-a381-8ae77300b5cc":["0","1"],"81c86cca-f827-4293-b568-ac62f7aacc46":[]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_6","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_7","pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_1"],"0000000000000001":["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_17","pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_5"],"0000000000000002":["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_2","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_20"],"0000000000000003":["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_4","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_3"],"0000000000000004":["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_3","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_5"],"0000000000000005":["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_1","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_6"],"0000000000000006":["pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_0","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_2"],"0000000000000008":["pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_0","pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_1","pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_0","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_9"],"0000000000000009":["pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_1","pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_1","pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_10"],"0000000000000007":["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_8","pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_0"],"0000000000000010":["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_18","pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_2"],"0000000000000011":["pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_1","pin-type-component_b21448dd-3ab4-402c-a381-8ae77300b5cc_1"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000004":"Net 4","0000000000000005":"Net 5","0000000000000006":"Net 6","0000000000000008":"Net 8","0000000000000009":"Net 9","0000000000000007":"Net 7","0000000000000010":"Net 10","0000000000000011":"Net 11"},"all_breadboard_info_list":[],"breadboard_info_list":[],"componentsData":[{"compProperties":{},"position":[853.049941,438.66969950000004],"typeId":"4690313a-502c-6ace-b9bb-d36c8b966d26","componentVersion":1,"instanceId":"aff8a528-b934-4625-84af-01f958e4a790","orientation":"up","circleData":[[782.5,380],[782.5,394.9638365],[782.5,409.92741800000005],[782.5,424.89125],[782.5,439.85482550000006],[782.5,454.81841000000003],[782.5,469.78224200000005],[782.5,484.745828],[797.5093645,380],[797.5093645,394.9638365],[797.5093645,409.92741800000005],[797.5093645,424.89125],[797.5093645,439.85482550000006],[797.5093645,454.81841000000003],[797.5093645,469.78224200000005],[797.5093645,484.745828],[917.5001605,484.745828],[917.5001605,469.78224200000005],[917.5001605,454.81841000000003],[917.5001605,439.85482550000006],[917.5001605,424.89125],[917.5001605,409.92741800000005],[917.5001605,394.9638365],[917.5001605,380],[902.509366,484.745828],[902.509366,469.78224200000005],[902.509366,454.81841000000003],[902.509366,439.85482550000006],[902.509366,424.89125],[902.509366,409.92741800000005],[902.509366,394.9638365],[902.509366,380]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[842.793625,151.64515850000012],"typeId":"afda042b-83c7-44df-952f-0baafaf4f876","componentVersion":1,"instanceId":"41fc28b8-a12b-46bf-af23-3da2617c8a06","orientation":"up","circleData":[[797.5,275],[812.5,275],[827.5,275],[842.5,275],[857.5,275],[872.5,275],[887.5,275]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Capacitance":{"version":2,"id":"Capacitance","label":"Capacitance","description":"","units":"F","type":"decimal","value":"0.000001","displayFormat":"input","showOnComp":true,"isVisibleToUser":true}},"position":[1165.012,254.87712039819695],"typeId":"2c229afa-5375-44c6-9069-3781267c16db","componentVersion":1,"instanceId":"07565f67-0738-4731-9f74-672de39f4e2e","orientation":"up","circleData":[[1157.5,305],[1172.5345,305]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"161","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Adafruit Industries","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[1075.654174,317.53555719008267],"typeId":"84ae97c1-8e69-5e6b-4fa6-dfe46d477633","componentVersion":1,"instanceId":"20642084-3e38-42a8-864e-12f237eae7bb","orientation":"up","circleData":[[1052.5,335],[1098.808348,335]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"10000","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Resistance","unit":"Ω","required":true,"validRange":[0,70000]},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true,"name":"Tolerance","required":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true,"name":"Number Of Bands","required":true}},"position":[1165,335],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"e95d33f2-d715-46ec-8052-7ee80f0ef8db","orientation":"up","circleData":[[1127.5,335],[1202.5,335]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1067.7176455,488.7010325000001],"typeId":"50189b42-5cab-48c9-8e0a-72db70fc6282","componentVersion":21,"instanceId":"c658a115-ed11-4c13-aea5-34348036d108","orientation":"up","circleData":[[1052.4999999999998,515],[1082.5000000000002,515],[1052.4999999999998,462.5000000000001],[1082.5000000000002,462.5000000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Backlight (GPIO3) for\nGC9D01","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[596.9049586776863,392.2291510142752],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"96dc7d5d-837f-47c8-b317-a9d24f1c8303","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"GC9A01","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[983.1596543951914,86.06386175807688],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"89c3afb5-35ce-4fba-a71b-117023af28ae","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"ESP32-S2 Mini","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1066.1280991735537,410.4500375657402],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"ede89323-f462-4ac4-a580-8d3a6368b911","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false}},"position":[584.2614505,394.9374995],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"b21448dd-3ab4-402c-a381-8ae77300b5cc","orientation":"up","circleData":[[557.5,395],[613.2041515,395]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"ESP32 PIN    TFT\n3.3V    vcc     3v3             red\nGND     gnd     ground          blue\n7       scl     scl             yellow\n11      sda     sda             green\n33      dc      data/command    orange\n12      cs      chipselect      white\n5       rst     reset           olive\n\nADC_3V 1\nADC_PIN 2\nADC_GND 4\n\nBUTTON1 16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1141.3685199098418,121.20735829938728],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"81c86cca-f827-4293-b568-ac62f7aacc46","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"8.77111","left":"523.90496","width":"741.46356","height":"541.38102","x":"523.90496","y":"8.77111"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_6\",\"endPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_7\",\"rawStartPinId\":\"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_6\",\"rawEndPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_7\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"887.5000000000_275.0000000000\\\",\\\"1007.5000000000_275.0000000000\\\",\\\"1007.5000000000_552.5000000000\\\",\\\"752.5000000000_552.5000000000\\\",\\\"752.5000000000_484.7458280000\\\",\\\"782.5000000000_484.7458280000\\\"]}\"}","{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_7\",\"endPinId\":\"pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_1\",\"rawStartPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_7\",\"rawEndPinId\":\"pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"782.5000000000_484.7458280000\\\",\\\"752.5000000000_484.7458280000\\\",\\\"752.5000000000_552.5000000000\\\",\\\"1082.5000000000_552.5000000000\\\",\\\"1082.5000000000_515.0000000000\\\"]}\"}","{\"color\":\"#0080ff\",\"startPinId\":\"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_5\",\"endPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_17\",\"rawStartPinId\":\"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_5\",\"rawEndPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_17\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"872.5000000000_275.0000000000\\\",\\\"872.5000000000_297.5000000000\\\",\\\"992.5000000000_297.5000000000\\\",\\\"992.5000000000_470.0000000000\\\",\\\"977.5000000000_470.0000000000\\\",\\\"977.5000000000_469.7822420000\\\",\\\"917.5001605000_469.7822420000\\\"]}\"}","{\"color\":\"#ff8000\",\"startPinId\":\"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_2\",\"endPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_20\",\"rawStartPinId\":\"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_2\",\"rawEndPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_20\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"827.5000000000_275.0000000000\\\",\\\"827.5000000000_312.5000000000\\\",\\\"977.5000000000_312.5000000000\\\",\\\"977.5000000000_424.8912500000\\\",\\\"917.5001605000_424.8912500000\\\"]}\"}","{\"color\":\"#FFE502\",\"startPinId\":\"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_4\",\"endPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_3\",\"rawStartPinId\":\"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_4\",\"rawEndPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"857.5000000000_275.0000000000\\\",\\\"857.5000000000_327.5000000000\\\",\\\"737.5000000000_327.5000000000\\\",\\\"737.5000000000_424.8912500000\\\",\\\"782.5000000000_424.8912500000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_3\",\"endPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_5\",\"rawStartPinId\":\"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_3\",\"rawEndPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"842.5000000000_275.0000000000\\\",\\\"842.5000000000_305.0000000000\\\",\\\"722.5000000000_305.0000000000\\\",\\\"722.5000000000_455.0000000000\\\",\\\"782.5000000000_455.0000000000\\\",\\\"782.5000000000_454.8184100000\\\"]}\"}","{\"color\":\"#ffffff\",\"startPinId\":\"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_1\",\"endPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_6\",\"rawStartPinId\":\"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_1\",\"rawEndPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"812.5000000000_275.0000000000\\\",\\\"812.5000000000_290.0000000000\\\",\\\"700.0000000000_290.0000000000\\\",\\\"700.0000000000_470.0000000000\\\",\\\"707.5000000000_470.0000000000\\\",\\\"707.5000000000_469.7822420000\\\",\\\"782.5000000000_469.7822420000\\\"]}\"}","{\"color\":\"#804040\",\"startPinId\":\"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_0\",\"endPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_2\",\"rawStartPinId\":\"pin-type-component_41fc28b8-a12b-46bf-af23-3da2617c8a06_0\",\"rawEndPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"797.5000000000_275.0000000000\\\",\\\"752.5000000000_275.0000000000\\\",\\\"752.5000000000_410.0000000000\\\",\\\"782.5000000000_410.0000000000\\\",\\\"782.5000000000_409.9274180000\\\"]}\"}","{\"color\":\"#c0c0c0\",\"startPinId\":\"pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_1\",\"endPinId\":\"pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_0\",\"rawStartPinId\":\"pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_1\",\"rawEndPinId\":\"pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1098.8083480000_335.0000000000\\\",\\\"1127.5000000000_335.0000000000\\\"]}\"}","{\"color\":\"#c0c0c0\",\"startPinId\":\"pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_0\",\"endPinId\":\"pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_0\",\"rawStartPinId\":\"pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_0\",\"rawEndPinId\":\"pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1157.5000000000_305.0000000000\\\",\\\"1157.5000000000_327.5000000000\\\",\\\"1127.5000000000_327.5000000000\\\",\\\"1127.5000000000_335.0000000000\\\"]}\"}","{\"color\":\"#c0c0c0\",\"startPinId\":\"pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_1\",\"endPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_9\",\"rawStartPinId\":\"pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_1\",\"rawEndPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_9\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1098.8083480000_335.0000000000\\\",\\\"1098.8083480000_357.5000000000\\\",\\\"820.0000000000_357.5000000000\\\",\\\"820.0000000000_394.9638365000\\\",\\\"797.5093645000_394.9638365000\\\"]}\"}","{\"color\":\"#c0c0c0\",\"startPinId\":\"pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_1\",\"endPinId\":\"pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_1\",\"rawStartPinId\":\"pin-type-component_07565f67-0738-4731-9f74-672de39f4e2e_1\",\"rawEndPinId\":\"pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1172.5345000000_305.0000000000\\\",\\\"1172.5345000000_312.5000000000\\\",\\\"1202.5000000000_312.5000000000\\\",\\\"1202.5000000000_335.0000000000\\\"]}\"}","{\"color\":\"#c0c0c0\",\"startPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_10\",\"endPinId\":\"pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_1\",\"rawStartPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_10\",\"rawEndPinId\":\"pin-type-component_e95d33f2-d715-46ec-8052-7ee80f0ef8db_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"797.5093645000_409.9274180000\\\",\\\"835.0000000000_409.9274180000\\\",\\\"835.0000000000_365.0000000000\\\",\\\"1217.5000000000_365.0000000000\\\",\\\"1217.5000000000_335.0000000000\\\",\\\"1202.5000000000_335.0000000000\\\"]}\"}","{\"color\":\"#c0c0c0\",\"startPinId\":\"pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_0\",\"endPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_8\",\"rawStartPinId\":\"pin-type-component_20642084-3e38-42a8-864e-12f237eae7bb_0\",\"rawEndPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_8\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1052.5000000000_335.0000000000\\\",\\\"1045.0000000000_335.0000000000\\\",\\\"1045.0000000000_350.0000000000\\\",\\\"805.0000000000_350.0000000000\\\",\\\"805.0000000000_380.0000000000\\\",\\\"797.5093645000_380.0000000000\\\"]}\"}","{\"color\":\"#00AE7E\",\"startPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_18\",\"endPinId\":\"pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_2\",\"rawStartPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_18\",\"rawEndPinId\":\"pin-type-component_c658a115-ed11-4c13-aea5-34348036d108_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"917.5001605000_454.8184100000\\\",\\\"1052.5000000000_454.8184100000\\\",\\\"1052.5000000000_462.5000000000\\\"]}\"}","{\"color\":\"#C28C9F\",\"startPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_1\",\"endPinId\":\"pin-type-component_b21448dd-3ab4-402c-a381-8ae77300b5cc_1\",\"rawStartPinId\":\"pin-type-component_aff8a528-b934-4625-84af-01f958e4a790_1\",\"rawEndPinId\":\"pin-type-component_b21448dd-3ab4-402c-a381-8ae77300b5cc_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"782.5000000000_394.9638365000\\\",\\\"707.5000000000_394.9638365000\\\",\\\"707.5000000000_395.0000000000\\\",\\\"613.2041515000_395.0000000000\\\"]}\"}"],"projectDescription":""}PK
     ���Z               jsons/PK
     ���Z71��8  �8     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Wemos S2 Mini","category":[],"userDefined":true,"id":"4690313a-502c-6ace-b9bb-d36c8b966d26","subtypeDescription":"","subtypePic":"1fa09ac9-b6db-4b4a-b77c-89392a61857d.png","pinInfo":{"numDisplayCols":"10.48541","numDisplayRows":"13.53099","pins":[{"uniquePinIdString":"0","positionMil":"53.93756,1067.68083","isAnchorPin":true,"label":"EN"},{"uniquePinIdString":"1","positionMil":"53.93756,967.92192","isAnchorPin":false,"label":"GPIO 3"},{"uniquePinIdString":"2","positionMil":"53.93756,868.16471","isAnchorPin":false,"label":"GPIO 5"},{"uniquePinIdString":"3","positionMil":"53.93756,768.40583","isAnchorPin":false,"label":"GPIO 7"},{"uniquePinIdString":"4","positionMil":"53.93756,668.64866","isAnchorPin":false,"label":"GPIO 9"},{"uniquePinIdString":"5","positionMil":"53.93756,568.89143","isAnchorPin":false,"label":"GPIO 11"},{"uniquePinIdString":"6","positionMil":"53.93756,469.13255","isAnchorPin":false,"label":"GPIO 12"},{"uniquePinIdString":"7","positionMil":"53.93756,369.37531","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"8","positionMil":"153.99999,1067.68083","isAnchorPin":false,"label":"GPIO 1"},{"uniquePinIdString":"9","positionMil":"153.99999,967.92192","isAnchorPin":false,"label":"GPIO 2"},{"uniquePinIdString":"10","positionMil":"153.99999,868.16471","isAnchorPin":false,"label":"GPIO 4"},{"uniquePinIdString":"11","positionMil":"153.99999,768.40583","isAnchorPin":false,"label":"GPIO 6"},{"uniquePinIdString":"12","positionMil":"153.99999,668.64866","isAnchorPin":false,"label":"GPIO 8"},{"uniquePinIdString":"13","positionMil":"153.99999,568.89143","isAnchorPin":false,"label":"GPIO 10"},{"uniquePinIdString":"14","positionMil":"153.99999,469.13255","isAnchorPin":false,"label":"GPIO 13"},{"uniquePinIdString":"15","positionMil":"153.99999,369.37531","isAnchorPin":false,"label":"GPIO 14"},{"uniquePinIdString":"16","positionMil":"953.93863,369.37531","isAnchorPin":false,"label":"VBUS"},{"uniquePinIdString":"17","positionMil":"953.93863,469.13255","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"18","positionMil":"953.93863,568.89143","isAnchorPin":false,"label":"GPIO 16"},{"uniquePinIdString":"19","positionMil":"953.93863,668.64866","isAnchorPin":false,"label":"GPIO 18"},{"uniquePinIdString":"20","positionMil":"953.93863,768.40583","isAnchorPin":false,"label":"GPIO 33"},{"uniquePinIdString":"21","positionMil":"953.93863,868.16471","isAnchorPin":false,"label":"GPIO 35"},{"uniquePinIdString":"22","positionMil":"953.93863,967.92192","isAnchorPin":false,"label":"GPIO 37"},{"uniquePinIdString":"23","positionMil":"953.93863,1067.68083","isAnchorPin":false,"label":"GPIO 39"},{"uniquePinIdString":"24","positionMil":"854.00000,369.37531","isAnchorPin":false,"label":"GPIO 15"},{"uniquePinIdString":"25","positionMil":"854.00000,469.13255","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"26","positionMil":"854.00000,568.89143","isAnchorPin":false,"label":"GPIO 17"},{"uniquePinIdString":"27","positionMil":"854.00000,668.64866","isAnchorPin":false,"label":"GPIO 21"},{"uniquePinIdString":"28","positionMil":"854.00000,768.40583","isAnchorPin":false,"label":"GPIO 34"},{"uniquePinIdString":"29","positionMil":"854.00000,868.16471","isAnchorPin":false,"label":"GPIO 36"},{"uniquePinIdString":"30","positionMil":"854.00000,967.92192","isAnchorPin":false,"label":"GPIO 38"},{"uniquePinIdString":"31","positionMil":"854.00000,1067.68083","isAnchorPin":false,"label":"GPIO 40"}],"pinType":"wired"},"properties":[],"iconPic":"c5aba2f5-4dea-4d75-9bc6-8c6f78bbb1f3.png","imageLocation":"local_cache","componentVersion":1},{"subtypeName":"GC9A01","category":["User Defined"],"id":"afda042b-83c7-44df-952f-0baafaf4f876","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"0755f9ac-cddf-41fa-8c34-4d71983a54be.png","iconPic":"2abdabbf-059f-44b6-b68f-d45f0cb3c7dc.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"14.96063","numDisplayRows":"17.71654","pins":[{"uniquePinIdString":"0","positionMil":"446.07400,63.46139","isAnchorPin":true,"label":"RST"},{"uniquePinIdString":"1","positionMil":"546.07400,63.46139","isAnchorPin":false,"label":"CS"},{"uniquePinIdString":"2","positionMil":"646.07400,63.46139","isAnchorPin":false,"label":"DC"},{"uniquePinIdString":"3","positionMil":"746.07400,63.46139","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"4","positionMil":"846.07400,63.46139","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"5","positionMil":"946.07400,63.46139","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"1046.07400,63.46139","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Ceramic Capacitor","subtypeDescription":"","id":"2c229afa-5375-44c6-9069-3781267c16db","subtypePic":"7c9bed20-c7d7-43dc-b689-820375f46db8.png","category":["Basic"],"userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"44.10000,0.00000","endPositionMil":"44.10000,-200.00000","isAnchorPin":true,"label":"pin0"},{"uniquePinIdString":"1","startPositionMil":"144.33000,0.00000","endPositionMil":"144.33000,-200.00000","isAnchorPin":false,"label":"pin1"}],"numDisplayCols":"1.88360","numDisplayRows":"2.48270","pinType":"movable"},"properties":[{"type":"double","name":"Capacitance","value":"0.0000001","unit":"F","showOnComp":true,"required":true}],"iconPic":"7ade412b-fa94-47ea-987a-d6c9baa14438.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Photocell (LDR)","category":["Input"],"id":"84ae97c1-8e69-5e6b-4fa6-dfe46d477633","subtypeDescription":"","subtypePic":"b63deb06-c33f-4ae3-8f73-25229955b1c1.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.58334,76.55539","endPositionMil":"14.58334,14.58330","isAnchorPin":true,"label":"pin 0"},{"uniquePinIdString":"1","startPositionMil":"323.30566,76.55539","endPositionMil":"323.30566,14.58330","isAnchorPin":false,"label":"pin 1"}],"numDisplayCols":"3.37889","numDisplayRows":"1.51833","pinType":"movable"},"userDefined":false,"properties":[{"type":"string","name":"mpn","value":"161","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Adafruit Industries","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"a5640015-ff5c-4848-bb8b-6d4b42e5489b.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Pushbutton (SIM TEST)","category":["User Defined"],"id":"50189b42-5cab-48c9-8e0a-72db70fc6282","componentVersion":21,"userDefined":true,"subtypeDescription":"","subtypePic":"4efcf596-32b1-4e3b-9735-2bd5fa764fde.png","iconPic":"a46afb92-29a7-4c70-92b4-1e1235f7410a.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"2.45180","numDisplayRows":"3.30020","pins":[{"uniquePinIdString":"0","positionMil":"21.13903,-10.31645","isAnchorPin":true,"label":"Pin 2 (in)"},{"uniquePinIdString":"1","positionMil":"221.13903,-10.31645","isAnchorPin":false,"label":"Pin 4 (out)"},{"uniquePinIdString":"2","positionMil":"21.13903,339.68355","isAnchorPin":false,"label":"Pin 1 (in)"},{"uniquePinIdString":"3","positionMil":"221.13903,339.68355","isAnchorPin":false,"label":"Pin 3 (out)"}],"pinType":"wired"},"properties":[],"propertiesV2":[],"hasSimulationCode":true,"simulationHtmlUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkitsimulation/136fd93d-482c-42ba-a365-5dad14a45bc7.html","simulationJsHooksUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkitsimulation/f9d4bf3f-59bf-469e-9f44-869dd8f99b47.ts","simulationJsonStateUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkitsimulation/2a1bf550-f602-49be-884e-a6bec1dae6c6.json","simulationLogicUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkitsimulation/8d30c2e4-c950-4b74-b8e7-566efa3b4ace.ts","simulationLogicBundleUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkitsimulation/c6573ec1-7f79-4fd5-aa54-a3173968a53e.js","simulationPackageJsonUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkitsimulation/245f325c-2c81-4253-8a7e-7d987b379c6b.json","simulationUIBundleUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkitsimulation/81067c30-2d93-4304-b1ff-a2a4c74fcddb.js","simulationSourceCodeManifestURL":"https://abacasstorageaccnt.blob.core.windows.net/cirkitsimulation/6402df8c-cbbb-4f80-94a0-c326ae044970.json","isSimulationCodeRunnable":true,"simulationRuntimeManifestURL":"https://abacasstorageaccnt.blob.core.windows.net/cirkitsimulation/ffd554ec-9038-45b5-9041-d8f2e3c5c866.json"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"}]}PK
     ���Z               images/PK
     ���Z�?.�� � /   images/1fa09ac9-b6db-4b4a-b77c-89392a61857d.png�PNG

   IHDR  u  ,   2T�   	pHYs  \F  \F�CA    IDATx��tW����ݝ������wֻ{fM�8����`��`al��	�-�s�j�V�B�����s�pc�q�9gl���ܒ�HHBz�U������s���W��~������@Ky�>2�;)+2TʌOt9��%�ⓜJ�䐗����.��Y�S�*9��H.���T��K�cJލ�\��9��`����a����$��F7_��ɡl���u.����_��o2�s�*Y�����8Z�����3]%"9�+%����?���>�Saz)xl	��R	a`�؀Mm ox�n>���!��ˡ<&9��]�xlɐ���Y�?�ѣ�}[0$��L�l�S)�_����T!c�`]Tf����J�*1K�S��r�s(JW��mu>��S�"9�ziH|�"g���w�h�n9�*t9bs\Ne�ˡ��w��H�k������!��A��֎Ԓ���H+�^>�ɨ`\��9�1��P�'�9�7Ո��RZ���Вm����t9��!?�r*{E�`�@��1�FH�9hw�w��Pg=���P��)��r(�K���b�Y�-;��K�W�	^$@�Pg@�κJ�H�@˵�S�Fr�ӥ��?���hh=Zΐ�.�R�r��~Y u�?�f"u��κ���ʗ�-Iʔ�-Є5o����S��L%B�e����� u��κ�q�'����Pdwf���7h)i���0�!/s9�oE��N�ۊ�YO�:�
P��W9�]�S��;4�z�= f:� ����� u��κ�%���]��@K�%2�u9���3�AP'��l�'@�u���IN�]�C���'�w[�T&��L a�:�f;	Pg=�+@��>�!A�� wh�jR�|�Z����A�����k��eS��8�������\�M��:��̡|(e�9�I�v��$򽢁ˌPwSQ�����M�/��M���/���n.����tCaPw�s[�c�w7 �̠_+Wdm�Ԗ�����r�@u�9�ΚKuS��|Vtz�0�X��s����>�򩥈��l���?��1�r9�c�6i��$��ÒC�^�1��	�u��
u0����}._*�1L��u�:�
P��9O?�S���W.��wь���F4o���:@��a�U4��zGqP"�>Nr*�R��������.��[4X��9Dꬱg�?aO��g �Þ:Kȡ�%eʇ�f4ڒ���.��p#3�����W�NP�98(�=uF�'i���K��!� +;�s(r�G�P�f�:@J�� ��}y#��$hI�Ň8%���h�2� u�:�`��� u"��-�
��`se*J�G� eF� u��P���D�?�)�rEvF�߉��A.���J�hp2� u�:�`��� u"���T^��2qsg��KM@hp2� u�:�`��� u�(5�PN�.h}4z0jn�Fb� u��P����!��C��2Q�2�\Ny�x㰆 u�:�`��� u&Rm������h�I��r�~��h��� u�:�`��� uf��TnX0$�iV"�\q9�բ�����D��P�ԙ�F��Tݑ�߹�ʍ��U�ԉ3@�P�31��岬��R�6iټY��KN�6�����D��P�ԙ[򫋳b�<�n�	���P6����P'� u�:@��쒜ʻRVd�h��e[xX�_]Ny��l� u��P���,v�*9*��lՂ�m^�p�"@�N4�� u�:@�e�P��u�B�9!9仅?T	P�f�:@�Pg%I��!���D�n�H�\���n��D��P��Y�ʶ�C�?�f#���HN�J�ю��D��P��YQ�C~��p�$�5�S.��g.e딍lS���_e�o��}��W��`_�-����;y�=s�6vG�f�ҽ��N(np���?���:�`��� u�W9Y�������;ؖuO�W�}�������f?|������){�w��7<�6��Ú�_��G����ף�G�2�~�Ŗ2�q�����'nzN7-�c_�௟��W0�N8��'D��f�:@�Pw�o�^��=ײm���~�q�&?�g���S�k�nc���H�¸�����2��Pv�
p|G��*�b_��&��::�k[�f-�
�8@"u�h��:���h�p�]�W���5���8Ikr�a�w7n<b����/�k�ةUl�叱����޳{���V6�٠���f&S7:2�r(_�r���+�f?}����{�CV?g���K��!R'�!&�[�Ãr�7�F��u � u�u���	5�fd� �������we��)��N��E�r�ϧ�f�T��S�Ȩ����)��� u�aP�C�.��nm����?���޹��ټY��5ɩ|�����+��L�\N�*��ȝg7�������D�o>���g���� u��P�ԥ'�і��o{��l�z��w���`�Q�i.�L�!m�5f��o�>u'�N���5�,�',�ZO�S��97#���e���3C������H��Nn�R�h9C��.���HC
W��z�=f�v��-B^,D����u�s�=u�S�.PW:�I]�2S۳{�z�V�1v��ʴ�tn�	�Ar*�0����sf;@�N4�� uX~M�H�O�(Q��������Sr(��u)1ɡ\a�!y�(R��QJ@]� ˯X~5��C���P����=e����W�4f�޴LL�r��7ژ贩%-Ne>;D��3�{�'�KO��d�T�
m����{�����2ҩI�C��r�_iLWGobVj?|��GU�R�C��:��:D��u�nx�Y����:͛�Cʊ�H�Fuӌ4����s�.f����u�:M��	��؏��aP��v��e�]ɬ��l~@�9�J�eX)S>�hczᾗ�U۪}6lLX~��h�IFX~�����^PG�ٿ|�kfŶg�V<�Q�y�ʂ;7oV���ʇFS�˙�m(�;�Pg��˯X~5�����W;B�퍛��ۋ�_�k.�^��a�&9��F�O�ì������q}����گf"u�u����o~bVo�ӗ�2�S�F4{��%9�=FS��+���s���',�b�U��OFX~� u�����a���
�(E��sw��לtH����5ɡl2ژ��h�&�iF�8��D;y@]�`�˯v�:���#)q��
��E~�V�&R���B�V<��_��ǀ:c>v�S�=uf�Pg'�����٩�Pz�ns#9�yvh�$�Qr*�mLT��N� ը��!R'f��_�'�K�{��ǘ��[Ͽ�'�}D�Q3�ޤ!J ���O3��ƹ�u|��C��,B��:;A���k]���H�v9�a�FT�rȟ�>�Kf�vW�^I{
�:D�D�L2B��zB���P>�\-yi���+��:���v˰js9�x*��t�ut�Ϙ^|@�\9��n;D��3��C��.Pg�������u�$�\�a�&e��F��RaL�OƎ�w�����D��e��u����؞��/�ΕC�.�P�VkD��2�5������˯X~3�˯��_�u�}�ٱ����ϗC.ΰR�fy/9�OSeL����ڂǕ�t��!R�H�Y��W,���(�e������9�/��S�U��s�Ҙn���ٵ��� � u~�Q&e��,D��u/��2�c�����3G̕a��ɩ��Jc��i3�k+�����
u�V}n�eu{uhP㼹4"f���Y>�ɨnvb���&��d�	�釷?��c���_�:��DF�foҐ��Tic�=̮MU���
u�";A]:	Pg�H�_����ؾ��{���!��l6ɡ<�j��Px+�kS��� u�aP�H����֛�S{�{�Z�F���P6e��IY��.�ґj�[���ٱ�޹����u�:@�N8l� u����~�ٱ��̻F�KqS�Y��kSt��)�̎��>5d���$�S�����jMa�՚˯����c�?c�ܕg��e����P>u��՜nvk�GP�? �{J�t�N�3 �؆��PW?g�c�X}��s'�����5ɩd� �.}��O�ݚQƄH�N���u:^��m��Y�|G��{�2���V>w�S��a�&9�;EB���cvkT�P�H"u�ԉdD�z��Ҥ�~�����ڮ�w���
S�0��fj�$�]r(;EB]�k��ڏ��dH�0"u�ԉv܈�!Rן Rg�H�������[^O���;��C�Y��)/	t$����٥=|�V��
P�\�:@��^{�HE�7���f��6tC�掶�e������������O0�������᠄x��� u��:һ�>`vh;w�R�	���Mfh���Jy�h�#%&5��}��������'D������`K/,���Aݬ���2�jf���`��g��]�����_����ж�{2�#��=2�/��.��/s���=�/U��u�����#u� 6 �3C���B}��7��m,��ڔϝۡ�k�T&׉��*?���9�>x�c��Կ�Dw!R�  a���c��ofVn�nxJ�8�B�.;#��$���h�;P_��Y�����+�@�P ��c���;y�Y����Y.�]$��P�se�ǈ�����`Vk)(G���+�9�6�=u����魖\5[�l�/nG�0aP'9�
� ן/l��A}���?"�K��Ş:8u�l %��÷��Ǭ�^����۟�4D	�:�CyB4�Lw4mfV�Z]6�9e��W,�j 5�,��k��?��B����X����"9�ۄ �7��{�S�E�dPO��3s�h�J�����P��� �R�o�G'�4]f��T<�Q8��r(_fdd�&�P'e�c�~�V�^z�Uf�F9���ޔ�9����u�@]�|N��
��;_23�_~�ɪg�	g�ʌK=�9Y��)����ۘ�ڞ�{�����P��� �R�w�'U�����Ծ��GV9}�pF�!�)�:�C�C��9�X߿�Sԥ�����5��P��C�� u"�bͲ��7>g��녳I�r(kRu�S�T��5h���<4�ڻ/~�
ƥ>Suw� up�:� �N�^���T�6�jO���uuqK~!�@wYV�O��]�*���/��8�͕w�%TD�P��C�� u"�-{R�#��돿M��D�Ie�4R���A��2I���P��+7*�5B'p	$E��K�:@:�6 �3ö�u��돾5����/쮖L�Sz����)�:ɩ��XG�\r{y��&+����j�2E��P��� �̔��2A����a���o��s.N�����\N�*�6B�S��Mw�WSM�۾��{�ԭa���X�a���ӟ u�:8t@l PgF�Nnb��=������@˧o}��f+k�`����d�P*Su�CyZ��AYͬꯇ�VnQa�����+�����{��g�_�sכ'q� �����`�:��"l�)�����W<Ξ�c��w��0��%?L G��e�]�fD�٥�$�rKʠ�2�0�} u�:8t@l P?��xRtv�a�?X(�9 ����u�@|�b�9p(ߥ�Ly���B��$>ȭ�:8t@l P_�4�����p�s;�sE����f��6pwC�mjXb���QyL�Jk�{�|��P'9d��B�:@:�6 ��ٚ����*�Jj��{� D "� "u𥊹��su.��R�@!@���)�`X~��y@r���C��o=PP��C�� u�:[�Cn4����
%5X~��+�@��+|�b�9�����C�C�.z���:@	�6�H"u���r��P��>P(�9@��: �6�H|�b�9x�p�s9�OL0PP��� �	l yꐧζ< 9�'�:�)%z�Prs�H"u� !l �:�R��s 9��u�G�� u�S(��D���K؊E�!�%ෙ�9p(/u.����`�H"u " l��6�2a֗��4�J��B�:D��;s 0� �l�
��T@���BI�"u�ԉv8� 6 �;���&��I1e��L���(��2�QrZp��? ԙ�A�]�:@*�
6`o�Z�.�0�ŧFX�`��|�����[���:/k�Y";�'E���e� u&xV�P'��@�� ���Qht�����ƃC�@j)����a�&�Ǻ u�'/������`���Gꂧ�Xc$������^V4+�\����JR�ԙ�!XA�:@�h�a`�	u9�eVqi��n��zE�|jP�x]IPg��`� up��*؀�m��P�Sa�H��f+�0d٨������ԉv8� 6�^Pa+Rs�&'��C�ρ�S�:<+P��CT��mf�:yR��^*�T�3w���pqPg��`� u��9���EN��U�^�@ץ:��"v�_�?+P��CT��mf�:�q��ON4�uWټ��yqR�:<+P��p �l��PGK��)<1X5{X��p?�� u&xV�P�
����DC�:p�hE���n�Rc�:<;B]��vy�O7%&��_oUL-dm���S.�#a`�+@�︘.��V5xYS���z��`a?k��'�W���˰�:<;B�9��`ֲ�PW��D��f��XtB���K���Z�C�q�#��ԙ�!XA�:�\s ����̴�%&�:�*��V� ��~����	Pg��`��L �؀�m@ԕ�׶���W�ô�361�.�r/��{ղe�}rԙ�!XA�:�\s ���(\[�WH������z��)�=	�3�C�� up& 
� l��6 �B���P��̧.��q�DvXS��e�ܗ u&xV�N���`v���9�PE"��?E�Z
�NǮ��2W�x�ܗ u&xV��@���D@�W��&ŧ{��n����T
Pg��`��p!�l 6`7�k+��OW0=�{(ʊZ>�S�4�:@�	���3P�`���TC��M-�=֘%+��G"[��C�:<+P'��a`�;A��(�;��YJ���7g�:@�	���3P�`���TC��t���k�qPW0�o_]�"@�p0� u�?�� 6 0��ꎗMu���­\�TY,����0�؀���s4ԭ�T"�%q��k�@�p0� up�p��� l�PG%�Vs���0�DM�A��98(��0X"RGG�����4��K�����D(�j��*�d�4&�N�G��`f�P��K>���އ��ɇ'!�0���`�H��.�9���u��DH����;SQ�T��E�W����}	)ML�� @�	�6 ������iQn�k)�a��T&�-V����	Pg��`��p!�l 6`7�������l�j)�Fْ�whT��n�o;�*;ǜ�$H�:<+Pg����m"��Tqi���' �v�1Q�z��U^�s�>QB#�3�C�� u�?�� 6 �#�FƸk�vii��|��\�A�ۺ�I���$s�����
��� (`�{ۀ(�#�z���u�꥝Q��)���=BV�F�����f�Z�L�?>� u&xV�N���`v����ڣuݵ������-�V�Xs������Bi0W7�L�� @�	�6 ����:R���&���;¼{��3�C�� u�?�� 6 �3���Yk"��Q?˜$\Pg��`��L �؀�m@4ԑ�R��4#FJ=ek?�� u&xV�N���`v�:RlbT��uz�ʒ���ωk�ԙ�!XA�:8 l 6`o0ԑ
������%a�s�JG�sSXd\��^buހ�.��ֻ�(��3e�n����� +�b��c��V�x���z����v����    IDAT����|����Ya<9�y��:�\s ���r�+,:!�J�Y�/�ZK����W�����VT{YS�Ϫ�Vt^X�M7PE嬈��D ]}�������N���y!������v���|��W�*W��3��ԤB�4ԑADO��Тu������S6�I�w|T=�MY����F�B��  	����5ͯ*�� +Ȯ�WET��i՘?�Ciu�ė�I)����*�����As�Q凶��� -�$�; ��0�̈
�Zӣ,+�C�{�q�?KB�M|JD�N�� �a,y�H��_,T�X����j����:�\��98��Yl�ԩ�&L���O�ޯ�Ν˪�4��.����iRI|T�����\u}�3�H���jON<hȬ���^�Q�L�����pg9��%ӥ�qԾ����i�utz�a����;���ԉ��B���'Lf#G�T5v�X@l.�޹��.xJ�5���5w&��*m�j)�����EK�.���FYK�����Q$���kk��h��Z��W�NK�"��J��j��ߐ�D ��X!1s ������ԑ�M�	�R�a�˲�ѱ~�B˾��@�)�W��}���
g*�2i�j���:����ѡ ZM��v0�H5���Y�'��%�B�}�	�:�\�\PW1k)�	���PGQ$#W��4
��폺�!�>�+���>�f��}�����`�
[0�F�����P�w�̖ʩ���*��:���scT�x)|�$@��.d�L9e�P7s�LW�g��5��6$��*���������cdu����V�hu����gFԭ[ :���u�~;��=j�mu� Ds_���@7T�/��D� u�?�P�� P{K���;�Q�������|��/�0K�������:��Xr=�
'#��%׃�̿��:�\P�{���T:����uE쌬�J�&�o��6yX쌈����v���^�ԣ��1¨(�*z|}Vht�xup&v
D��?�PG��D�����cX>Y�r$z|�hE�����,ut
$U�lxE����G�yRuʕW�ʼ�28���P'�@⡎���.�՟h9�������AW��ii�?`��C]�� }�d�~˰��D��~B@��.�N�3�C�a��3�~�^�7K�7�r��ʟ�6�ŧF�>L�]�#{�#��2�\eE�0����؋3B��=|A�
��'9�29��^�`�{%{������}�::�1j{��a_���K��;7���meź��������ӱ� ��?H�$fE��GkW�ؖM��;o��~��k�X�����;�������m74$�,�{�>��r�%�$\�$��I�ݾ�OKy���)���F^)��H�������2KBE�4'n���E�wt��S^������������.G|Iht�d*SP�X=�tͅZ��y`���wl0�^�;nj�<�)�.���m P'�@��@U��*���5�>����엟�?����-��j�G<iN�������uS'�}�=$67��Ŀ��ҡ��#Q�	�oZ���O�SA]쌨fr�N����}d�w��7��{)+�(�(ءe=�=����P�x�Za￳�񶎎����h��QT[��.�mm P'�@��lN�&tM��>��Mn�o�^5�|�^%����Yh�B�%9)����`x���=\^F%дܳ���g�d�C��t��c?�����Mʔ�)</�K�D�OM�5�\�t_|�>K����qM`WqQ!>�p<��@��g ���f�?Ȱ�=ξ������ܯ	t�TX2�WKQ��J/���匝��7ʂ�y�}Z�9-j-��.�� ��6{(B�!9��I�/S9���`�$��C�Y��㻧WS�����c�rUs<d�����/d�F�ޯ1'��E�G���ws�}��:�.�^���Xx�b�c�C�:�� 3�q�lu3���|��}��;��#ڇ��jr��_�<��BG|<%��=$vj2��*/֒���|��:*��=�EA&9��}��[V��>0�5L��;�G6�gz�}{���Up��R/�G�{	��/�_��H�/�>ց���)���
�ԉ��9(�.��GO?~�n�h���l���K���>�D�ô�㓜�b=x#oD���|����g-��Mv����<G�>��'��z��ּ��	���ã�%C,�0�}����ez6:��m�������6�:@�������Ÿ��U��l׮�u�G����?
hLF\�
j9���`���9�$�w�"����z?_8�:'�$�ҳ��ar>�?O?�h����>p�Z�w��'�//��G�����i�ĉl	�k��K��u M?�ܔ�Ŭsg�B�N�3���AK_���o���ٽ�]��/���toM[:�*9����1r;���&��Q���)�#R�|���\|h���੼��j)�;���k�2#ڣ^�Տ�<���s�=�M�>�pE]q�cH�]�0%s��8O�X��N�3�����>����W�G��j��G���Mhɖ�N��'4:�s�!�?���C�[_�xv�:P���o���G�5��E�B_���V�fM�������՗�����H��^@���P��>B��S+�I�ک��kW{�Y���������&s�sgɏ����W:/���/�Xꈜyj�ѩ)Sy؈�*S#M�	Xް+U�0��/.;�����"u��_(�s@�Gy�j�hE����1�tT)��(��R��怺,����zh?�mF�U�~��/����/�qj��r+z7���3��B@�_��:s�LW��"�	on:�ڻom��K���|��Aݲ2/��r#x�pF�=��T�ր:O���Β�6����o��xh�����޽Ӑ���w_��%��:����\`���v�8a��4-cǎ=�>�.��U�Z*��!�A�6���ԭ]4,���+Oq�����^���s��5u��F�F�����i�,u+j���R�ˌ�����O:�������s4⃺���А�h�q�ci��5`u��T@�ܹsY՜f��a����
�鵺�3[���G�B~��B<� �ۖ�s�wH���=L�y�@���ĩ��k?3�c�|�QJ/�v��I�;���-��D��Z�Տ:�bjG���Ŀ����`y%��}����Gw���Տ��Cڂ*���bgD;r�������i.���@mx���&9��z�3�h;o�2��_yS�����v����]Η���Bs�s�sXnn�~]4�b6g�Ik��E=�n"P.|�)��������2�/��w�C涉�jʨsظq���:��J�4�|u_)�w��ߚV_J�.����e��rXO���n���`뿚ꈸyG��^��(G]����I�k�h]4��L�����K����}(�R�-��-m xv>��	�ʙ`��~U8��叭2��ײ�m��sP1�I���U5K�+|}�s�--��=#��З(�,o,�{ž�2�Ӄ7\��ɔ���M�w��*JO�;�B"ږ2�ۓ�[G{�����l���*��'���YG�>Tw���Z���+�|jN#� s`g�����y睐�spe�z��֬J�Hp����X��j�}�9�����`��K�'�E&��u(+��C��+�>��|��~uU��j�]2W-�U�L�r�����XR�K�~:u��
k���sOޕ��o�>v��V�{7�}���� u� -����GWpgd�k���=��-��r߻|���t���eƻՊ�?-¤!�;	��M����	�efR�E!kA���h�2lg�U��24��'�����v)2N�~�.���[r���$�n/{辫4���b���� u�:v���[��Z�M��ݽ���䏂�j�������M��/��r�%�����>��Z:�e��d�A-I�%���Q�w��;3~�`��xH�q�c�Oi�Б�ʽ̥q�K��7ۥ����]e��\��آ�~˫��*��C�1�:@��KL�_��;/{� ����_�[���tO�����%EO�_�U��a��!&9c���d�7���i�����i㍥���k*�#���D!Myrx�+K��匟��J�����M�t��s�|{�P���*��.�&-ʈ��7\]��J�e�S�/<��]����X��/��;;s�6 �ԉ��&E�?ڸ�����K�����ٳ[��μ�]�)ɭ�um��M)r�����=�ʕn�2M���?w�˲���ﱱ)�oiP��|Mu�Qڢu`����l��ȏ�3"��#?�	[� �e-����}ji3=�N= ��x׭��-�׳W�?�>|���������^|�A��v5xR�Y�c��9Hw��뮻�A���i�=y"b��am{���ث/?�>|�U��m{n���zy�v�"���=�z�_�L�Ѻ��<�U+=LS��{�ؤ�/�9!��K���}�G����:R����B*D���Au�B����Y<�LD;{(=��`P��s�A��C=��h{y��Z=J�"���O�A����B�����򎐹�h�JZk�|��=����/�N����c uɁ+�.9����Zs�_-�^�︘����)�`j�Z�H�99ٰ�ޢ$�z)<6��2�ޢ3T�P'��C�3�:@�H���}�H�۠�ֲ2�9���LI~�]g�a�0�>PGJd�W]0Jt�"t��a_=�L%�����"R'��C�1�:@�h�#�]2��������MF�Tk7HT��"�Z�aj�3�DSĐ�?iP���YͽO� ��;{(=� P�3���|3�o_��QW����
�ј��]� R29�LudX"A�&8vF
��(s�����Ӏ:��J�9 ��� u]�#� ߊ:��	v�.����@��顮KE3�lU��صQ*��\��cI&����%ݖ\���g泼��,g��]:s1�_�8�J�o�g�>s �ԙ�~��H��o�CG	R�{)��VR<��b��x-u$�ee�9�R����#�ٔ9XO��E�S1^J��9�x�	�O��N=����>}�A�_!����P�.9)��?ѭ���ғ�tQ��$-<��£��.R%@��lPG�%P
t����;1XE�GS����d���鷥��D�AJ/%�@�?��ꝇ.��f)�dnH]5*:Gy��4���G^�F����O����G؉'��Fi֬Y,���M�:@����3\fju�V�(hK����(�p�s_�AQ�ք/�򖇺.yFȬ|AH��̕���_9���:�O�Z����O����L�u���A]�İ���M�:@�Y��K�cc�^;��+�J�,ZD�Jz�w��V��kXk���O�$]?�VP�%
Y�1P9^�<l�)�¬f5��~)�Q�Ky�KǤ)yct�x���qE�������N	�M�<��'����n���u]�;\V�7F�܀Gy_��;B 7��Ƒ��i����)��1Q��_iu.UҺ?M:�Lk=��~�jr�IZ�"�yc�ĦB9C�@h��<p��/�B����o:Aݜ/�:�dEx��K�_̦M��E'�
����Y�z��a�E�Pc��_�o��:���!�a~�sΥ���եS�/K��}��'��K.�S"�w|�V mu�qs ����_R: ��%yJ����M�:@��RL1�:<+P��� �~ԥ�$D��?+P���D��:Ѿ�er�L�� @�P�l�:@�h_�2� u&xV�P�ԉ6@�N�/t�\�:<+P���D�P'��L.@�	���� u��P��]&���
�Y��.l`�e-�U��1�T�.j,m����S2��i	�;>��?!��&��+��r���C�JX޸���������{�f�X��$��.o��.�w	�?o>�=k6�q�v���UE�q�R����.@��IL�uvԜ�/d���3�8㠹��Ν�*�4s��yg,���'M�4p�_y�acԙ�Sc�=ǣjɹ�,>��_.(c��jz���=*��u�Y���D�a���k]�:���DB�đg�wzcǎ��f��p��?�S u&XFuSGOg�ƍ�/�mP'ޯ�Q�ԉV�P�C�.�����:�~͎� u����� u��͎P�w�µ��{�ϰw˯�}�P��$d*�s��|��Xन���G���nʕ���ƛw�NˇmΉ�����|��.�aO��:�ĩ�v�3g�d���jҞ��\˯~�QbO���nΜ9�lfcJ�����=TayG�?�Y�X��=ܾ�7g��<�xc,pb�xs3^�D��#c�hf��z�5�c��<����V�{Ys��U-
��Y�gQ��c�3¬&/�Z����k.���A�a�#���:@����ԙ)Rg�	;A�LѬ0��Xk�������󲦸�U,2�̈e-����xv���lY���7��k��I�K�L�I	�ZꈄɐZ���������W'��]���`������*�j/_}���P<��� u�ԉ^Zԙ�h%(�f-�$��R�
��3��mr�K��9a�Z��<�U�^55����:��ҋ�*�k��>D>�f�͸��^b+j=������g�5^@�P�l�:�PGѵ��AuHO�R�c
L�s��V�(Ҷ�A_�h��������rPG��ID���1?�nL�x'EX[�����~u��N۞����P�IaO]��h`����j�Q`E����!�W�����(��=��~����=FN?���I�FN�aRZ�eP�/��6�t�ԝ?�b.�k���g�P�ԉ�SG�E5����#�Ƨ�����7ڟ�2ި�2�H�@��i.��l����I�T�bMj�\�r��k����*:
�H]��{lLݚ$��/�|;��x���C�Ǻ�٣n��=���`�]uހzd9EaX:=$r��� sg���C���	N��da�U?���FowH5��V�T������rQr kj���&ɜ4�S���O�҆LQ�����"�S�n�����s�U5P�Q,����?�ԙ!��w�l�~�A����@G���W�d����:��Z��Oe���'�6)b���NG���-e�3���8�0yb�A[!��v��!R�H]�.g���?탺+1�8�K'zE�� ʻk+�#R=�}�y�&�y�|AȔ�U�٥�A�@�P�:��v�珚<,2Θ�n���t�]�a�Sb��:J�'zB��g�t�
9-������5^�{��3ؤ� u�:@]j�N��w�S[�O�"���	W{?��X���Mu��cY�W��$Rm)�6��٬�FF���^��h��*a7o�f׮-bkZ���UK��:�M:P��u��
t;�vy�]O�h}�pE!ko�n,V�zuKò�x�اΡ^��eg�A�JKfhcg����\ʌ]-9�R�C���rY�py}tB�+�t�Lvh
ӱg=���&3^zY�������}�{۳g7���7�c]�֮Hby��a�	w�P���P�3��.J.JG��M웯>a�u��G�w��{�mٴN@h��K=�3B�K�1�ok�����I�\e��)����P*��o�M
�P���`D�B�iI����Q�8p,e�+3>&##�7}�%�������}�Z�nX��&mT���͙�+���d���e�i���#{���[�w�P���P�3��1jz-��UQ����{�k?��-{�����%�O��R�Z���V�xY�9�%Ny�th�	��Ob|��]��پ�嗨r�����3�Q�U-^V�e����!�\�r��(Sÿ�sCd�����B�2��,���{������5�:i����r��J�9 �� u�B]�M��u����/_�����%����5����ؗK����)S�)�ګe-vo����!�O����t���QZ���#O�|�%<���q���;���oX2��_e���O�Z�/ܹC�9�:@��X�k-�ߢs�
�� �    IDATu(���ϳ5����$ˈ��7~��Q��פL�P-�A����?k�oGu�-u�'��� D����%N�d�G�����.�In��5���/�ؗ���h/o{�ۨ��ܡ��@�ήP�{���>���:�����u�
N/c�����ʕa�ݷ_�⏞{�nnDA���*e��oE��y��~�;T�J�7܎�Y�;x�O{�,uD�Z֙%�"��Gw��k����`�������噭w0�Z��ƥ|}h�0�v�N:j��)�v�s��a�3����������rʀUDj�+*J�WE	��Q.��LT�ns�s�������۷W]����:��*O���;ނia&e�����������WyU>�4PǛ|�6t���F��#������Zk2D�S7W���]�~fz�O>|�۰Kf��h�IGMy֠�ܹsY�fC��Y^i�Xu�:�m�LP���\�����ݻGWD��y���伤�<��O`���:���E�����w�������Pk����Ow���V��.:/���t�>x-3��pu)W?��N<ण uX~�u����]5�[��v���gGR���U,��'o������d	��EFO�,+�'=���?�r�Z��»�߆�>��"3�m}�f�~�{c�<�~s �넺��`��nKE������\�d���_p	[r���H������~����G�}�!������G��g*�~|��N���}d�wz�{�||�߯{"b�@/�zF�o�ׂ���y�Q��m�&o>��ڐ��W�����HD����o�3e�,�j�yn�YI�*Z\�
&�9��Y��iH���fI�����B�_!�s�u3ϘͦL��j	�A�p�Z���2���;�G�{��/TH���ҡL޽���F�F�E��<})_��e*|%5�=,'S�lD_��/�L2-k�:ޓ���.�#o���׹���	X�a��s �3ԅ�(b�iQUy#,<��_E'�0e�x�Ѣ�i|�^cF��_�T���?H\N�*3���X�(�/9��F�U�y��/�~��,|yj��J���>��->�+ ԙU���ag�<{�&�<��uⴤ5��sz����5�L�3ԥ���ʹ| �{3����6���z����8>���a.����(��:�Y�ԑ�x�3\yވ���	��ӏ:��Ho�ٝ;w�����\�h���jV-\���):������jg!R�K��ɣ�"uT���Ø ë/?���w��+m����mF�F�������o�[^�9�Q���Jg�դ��?�\ܙ���9k�~��;��D/<���K�Q�N�{ u��@�.�6ǻ�{��؞|��k���9W�<�st���[��*�A˩<�(��BPפ�AN�����O׳��陪D���d���&Kc|�!�2��skW?j�(���7m3f��:g�4<�xr=[Z�<u�`���\[9_���^�j�?�xmW?�fi�m�|A��Y��u���pY)_?
�	[�(��[TW�͋���[y�(�����%���W�����=�|\�_���f����y&��C�-X(|�� 6��4E�*:ݵ�Ew��ןr����-�?��.I�P*��ȸ�����Z�
g�툌�tP�=��xH�q���y�ՖѺ`:�x��e]_�������� u���s�@��8�/���t�G[6���C�����{Ie�B���ݙ3������)O�C<}X�tpeIMuZ
���{X�C��L���ShT��(ݲ2�&�"���۬I���2�g�.]^�o��T���s���~���9@����6����)��G�^_�[�-�3��իa�N����篽N[��L��DF��M�����i���|$��*Hy�։����;�Q�-��n����>B���_�tz�]�~a7��M8�aN��NP'�@�K����le-�?z�эI��;~`׮-�w��It��0����j���뵲�7��{�q��+���]|~�ZPG�	�(�|A�����ެ���-��w�|O�·��K�S�-�v�J~h��[n�|�|�Ο�75i�/���� u����m�.�����S�$����pOq{=�������N�������w|�)-�ZE�Y�h�]k�h���7"��4$>s]���??|Z�#-�ARs���o��!����ҽ��`;~����=7\]��~m�~&�Zgbbg�H��g a�j��K�S}t��{�d;�˥�ɇo�Wj�e�H���F�/�v��d�#�ݙ��Yt9�b#_/��������TPG�v���:0I`����v�)�K��9�Pr�D�{�S9Ir(E�Q�7�s�2�S�z�Z ]�2ʞ{�����>V7���Y讒Yq�P�{ 0����U����f��/?\�|��j�$���z��@5F��ҵ��*��Z-�p�iɩ�\�X�/G[��C��ǕC'fçE?�ӳZ�3�S���:�����~5{�Rٯ�y�<6��եN����g�Q���J�q1��Q�q�ִ���76���ld�_x����q��z��kٍ���K-	��������������5k�1cF�:��z�]���B�؀�6�_��@]��gw�ܬfWؾm��^x�~�e�zv�U�2���u)<&�9:���T*�a��n�qAHP��'�����Mu��y�--2��X}~%t�D�^�T)2.ʂ�b?�ٝH�yKYͼe�U4��EƗ&��)�=�nEv��B�؀�6�7��U,4��m������su��`Q���l}��\,Z6�B���;���x�ɬ�Ȝ��&�P'
'
�����Y[yr�GF��az�_ϑ���*zl�}�d�SB)02�]��hx�Qh���k�ye��\�M��';ԉ��B�� l�h���}��h�۠t�u5��FN�&��ܮ�hIW�xMu$:���a=E����Ay%O��ư�%H����@��ԑ�E��o�������hc�/�=��_E+��Gj�����|�hâS�����Gw��a��[�e�Sz�P'��a`��TA)�6G��xc��L���(�t����T�9',,b����'�1s �O�����{,��@����`5��Х
�D��DVZ����2PG��4+jS�Ǯ)�g�Afq�[�q�Bc�B�j���������0��@���$��TV+Q�S�Q��.ŧDR���>�׼�jI�#yGȬ1����͝�l�ڔ9X�����䈃E)��;��� ��L ��@zB]WNե��Y����#cj����6z�<�n�r�Z
�S4�;1���P�<8Ɋ��U4^��k��N����`f�:���Z�j 5��*L�����ٹ�ߨU�:��ǁĴ�:ո�V0#�K��̑1Q�]�Fԏr�*�`ZX��}�_��KG�~����� 2`�����wX�^;��?j�\z������eV<;��*��:o@McD_-u�Eu�h�����⥨��Ivcb�S��R��ή��&P-�Y u�?�� 6 0�u��Q�%J��Z��Zr����g���o&�w����A.���y8"6z��-�����I��i�EA~��_R�q�Q��+��ՕwD��/��9ae�Ó���@���x���}�T43��.����G�dn�ŧFX�ԘZEI���C�1�g�̰���_yc~����[�h{�����-�Ad� ��p!�l 6`f���s �3�C�� up& 
� l��6 ��k]�:�ԉ��B�� l P'��L,D�L�� @�	�6 �� R'�׺ u�'1����0�� �N�?t�X�ԙ�!XA�:8 l 6`o@�N��u��Ob:P'��a`�@�x�2��3�C�� up& 
� l��6�H�x_�ԉ��t�N���`�:���eb!Rg��`��L �؀�m �:���?�� @��.�9�� u�����B���
��� (`�{� "u�}�P�{�C�?!���M�2er�EO����(�G!���=���_�ԙ�c	a`��t���#�EXlb���N���(�m?���R������2y��=*��E�.g���3#�ba�����&ko�_��li��J.���%����� k)x�+<l��g��Xxt��3��H��.�9���u9�e��aU��5�c����z/k��Y��0�b=��;\a�)V�$�ZK���u^���Ĝ�l�x-u�k��&�`�:���z�	�;�ܿ"(W�(�V�&9�2/K\b�G~��:8 l 6`o��:�*WP$�Z�}�xvH�C�>��>����	$=ޖ"?+�6l���:�q1V�	���W+뼬�"������5`�V:/���Р�-���0�� l@,�Q0���g���G5^V2'��D����8)�B~]��N�j�
��],}�.SQ#L�����V�c��#�6Ei����V�Խx�:8L8L� l }m�`PG{�(�j���dE+g�?\�����!݃)��%�S�E��цCZ�6rr��~�T\TY�A��x�up0U.��+	�:�\s ���t]��i{H�ҋ֨�V~v���P�=FfMJ����Q,��N-�����f��ǟWiu�\^el��?5F�Z��S��1�V)h�Q?��co!�N�����g^��j��ܢ�[�ek�֦7ԅFEեQ���P#f����Ӣ�V,��$H2=ԑA%{"Y5��$#:��V�XI�%�Ȟ�ԉ��C�؀�l��PGˠ�HV��!U��)تF����=l	u��E4�t�I��� ˫��o���Eԉ��C�؀�l�f�r�:o���m�����o���货h��bf�
Jof������bMu��'��jr�-yR��c�.:a��ч0��@*l���M`���22ÄYH�l~�>PG�q�|�ڗ
�bTj�3�wf�x��SX�`i u���X���K���JA�1h%N����8,B�������#�'�?Qz����+S�;^JC�:�\s H/�[���gw�=ȶ\�${캧T�PWt^X���O�x�s�~�dE��D���Q���(�頎�]))_�0��aͅ~um��`��pY�>4^��o6�0Y����/�7T���\���
v�m+��W��3^�Pg�<�9���T�Xƾ��۔������mv�u���;�Ut��m�ڵź�#�b���� �y`W5z���¨�Fد��c�����PG�M�!�ٛ;<���Pd�S�x�S�D�+eʊ���֢١}�^�T}�#R��d�q�MM��7�g�w���߱�{�}ۖ��`r�����s��\Ϛ/]�_wn(?P�����xR}�kJ�[��[�sZ{\SvNc��[z���X���s����&���5�א
�����jfs�k��k�_5�[z\W>}i�k�?��i����Q�kK&7����sAόw���ٴ����*:��}��w)?�Z�09�{�m��{o������g�~�����l������Q�Z����@Rˣu~?��ٝ;L�Gr*!ɡ\ 9��n�2�吋#c/$.u�H"pC*��gI����ֺ�m^���r*�����?�C"�����*��Ӛ��<Y��Ӵ+4��^���}y�/��}�؋�?Ȯhj���HH��J�9X�m���zjӃ}^�ܖ�{\�����ߺ��ߺ��^�<x��=�Y_����m��h��Z��u͆�k{\�y����)<���5$���m��=��}�-}��޵w������z]s�5w�������ti뽛{\�&���5Oo~��5����t���9�O��{޻tmE�9��ǜ�Y���ݻ~��6�y�]��5^���>���3>�\s����K�'�9h�w�n�ܓw�+LZ�W�N��RBe&��jC�����J��)���xc������������ք��a�yl򎊽'e�#x��"�l��Ċ��(�1��i����vC���������uk�~�L,����s u�� �Kݳ�����չ}���[՗���=���]�~��>��uv��(�=)s`.U^�]�����";xxC?=6)����)��6W���NK��|j�K�e����o���C��o���;�˚�Q�R1�=i���]}/��}��'��U1�{�,���A�9���y ԥ�����޹c�OM�=����"������ݓ�?��w����+H��3M)��~�o�=2�/ZxCʊ�L�|�e�0~v�ZP�9ZV�A<���2�cb_H����/�Q0$>5��$��H�F�w����_4?��5ӣ��֋�F�V����s u�� �K][t���޳{�������Y���_��y������'��OiW��_J����ʽ�O���C�?&����W��eԖ/�@]\CZ"u�C9W�>��'
�?��k-&��?^:�g�t���6{Y|\���~s ��@]z�����ӷ7�o��*�p���^NGoԡ���G�����[�bgD:���z��;S	4���K��z��:��E͕^�Ί=�c7>-�"��>][2��|�����'�>�}��G܆]:�H�J�9 �u��.}��5[����_v�勯6�^�A� �ה���]��G����c�e��Tgܫre�^��}d�wʔ�'������f���$�S�ֹ����ֶ���3�'���h�O?�b_��}:
P�9���P�YM���M��o~���~��7Uл��5zן��oY�/��³��Fܹ�
�k�%|~�hf�-�'o���
�!��T�0�Q�gp�q�]Z7+���hrł�^�~T-�v��7Oއ�b�K��3O��ՏL�J�9 �u��.=t��Z��t-���<~���?`F�G�����5V�T����GF�Hd$~�'o�U�j���;%sCց:��8yG�/�ׂᏵ������g�O��Ѿ�~4�"�?xP����s u�5��A�<����i������mW_�$��yG(\� 6qe���%�vrA��@�3����]N�#�*O�<��*?���~)xYG�>C^�O>|�k�[�X��*��)e�I��h���g����gy��u���>�֪�Ip7o�u�7�L�{M�U}�o��Gz\�����u�W�L�{��Q���J>\9���u�����5����g���֞�����u�}����k��w��޷�gb���^�<��=?GW��w��3|rS�y�҆��sv�u��L���'�pB=[��A�x�?��Y-3���o���/�y�A���{���P���������::��{�Tr�w�W��\P�:w��ګ��ԮFY���� P'��o�ę$I����gŅ'�l��g�Yՠ�����U�㚭���������W-��~۞�	uUe��Y��f��^�x��^PWWz]wㆫz\sӵ��ٯ;n�	�ֶ����[o�q�UkV�;��?xo��K�{]���{n}M������?�P�y�ҕk�3MZ��^�Mʸr>�kW�Q�7_`F��Q�W^���r��Q43���uoͳ�ʹ��9B~Ɉ�L�eT^m˯�Ɏ��S�DX~�NG�+�W�U��گ�+Z�����u��uMaA��5����������5e%�}ޏ���ur,�뚊��״.m�uMNNN�kH����u�ݯ������_�ldu�������_����ڢ��^״�X����0�缯^��3$U�����/�����.�Ri�}�����ңLo���*sWspg*w��B?����RA�r΂��1�_������wH���{��j	�Q�x�YS9#����GC *��:s`W�[麆������u��-?�y���JKVsU���cC�����Տ����Vyk����?��gz�F�Ђ����;(Qz�U��9�4���C��g?)EJs>gJ�lm��hٖ�>�l�Ð�����Q�)MD;�P3���������VnQ��������Z��V�d��M�g���R�~̈�$�D��0�+�pWs9�AެT��2PW������6    IDAT�衸�껯.xj�	�>�b�U�B��R��}��=,�ݷ����x�Q�m��Ɛ�9 ԙ b @� ���0_����0�Հ�����4&��KA'�SY�kdgd��<)��x��Ĭu����fŧF��2I�>JC�)��|�j����L���h���Y�Y���k���?�L8,@և�%K�@��l�J���Y���\��٦�[�����~%U]����g������Vp�����{I%s�˄�O��[<4v���*/�]���*�*�{̘D��ܣ��/ˊ�)��I�C���� ���-E>ME�ͷY��nM\���L��tm�~�@��P�h�"6}�ts`�dgg[�̠��J����W��ݻv
9�GZ*kK'F��b��kI��{�����'��-pL��{�M?����HT_�w��7�j�j�腇E��?2�܊j>�!�^�m?]���|�N�scK҉����r�_f�.E���� � ���P���ʧV����h�]k�Ρ��ן��V�C����2�g��`�;S�I)��ޠ Tpt�:Q�{��s�փ���|E���?�r�Ƕ�:
���kqV�ρ����4�%�	�oL�3�C��{o_���ޥ����/����Q���R� Yg u�:@������{�W}�����5����C�]���Ֆ��/?b�//�'�^�ծd�/���2ު%AZ}ܝ�/ސ2�᱑�y뽪�]�a�G�փ:���`��B��Dw��r�@�N��I��;SV��	�̛/�K�����=\��Wץ��U�/>{����`o����_D����Cd�9 �� u|�_�hZ�ׂ�˸S}t�����7_}2xo�ѡ�[�\[ �Nc~��� s׀���=!���P��#�;o���ѕ����!8�r�j���k*��gmY��&�����ȏK2c�$�<�팟�3$v��ۡ�w�>>5��7uɁ���v��@�����{(��-�_g���̚�~����߼�7��$A�Ј$ADx "�� *XU�]9�[��s�MgrDQ��	0�gŀ�"��_�b񺺫���P�ޮ}���y�^���S����}���%{+m�؃k��=u�8q�8|��e���E�����	$c�AAA�<���_����C���_�_㗒g��"���Z�'���X
"D��?
���wm.���C�e��#l3&wm�V�j����q"^gNL@�0�.��
�f��̙�>��+�G�߸Pg�@`nvM-�6�/+�J�MN��RS�ߖ����dK��1�o�Ã�6�ӻo�g��.=\;����&��V�����!�d�9 �#�#��u�~P���o<S�8Qr�gKY�J}&��1��wo9�0����o�i�c�.�/���15�٠�鄲eN��F���#�J�f��Py��5K���9aE�v������t IFAAA]��b^3<�z|��Q�[�~�=<�j�.j�����#��G��o�M�ݪ��-Z,?:١�Z+m�e�t	uX��C�'4��d���4��R��mI(R���&�:�:�:�g�~�Jx|�3R�.��͇����OA��6͠.��J�'i%L.T��f�r%�m눢���t	u(�0��R5.�`�C����rR��T������$�������N���p�jxr�s�×?F����]-O@�5-�B���#�Ъ�1(5��ߴ�(�h��$��Tf��W^�P�r�󫲿����q�˕k�~Vc���t���IFAAA�:���}j����ׇ���|4�>ۑB)ԡ0P�3�j�>`��="^�/��r�C�N�e������D����/�a;�j����M�A{-��Tl۰�s�u�!�h"�#�#�S��ƖB��u�g�>��@��BjAJ��]�DՀ����_lW���P�2˷W�P�¦��B����5��չ�	��� �ڣu$��IFAAA��������:)�2��m	��i�C�U�4/�e�ǡ8"i�Ca�i�3Vd`���.����$�J��Y�!��$�(wr%��^S��WB[S��S�W<]�	�{}q�ݰ*6r޺���Vx��I����G�ξ�/�K;V��GX.c �������J��0IE��u(��[]��G�n\�_5�re�w�p�����X0gN������EE3k���ƭ�wm!�#���Ք�3�����?o(<+�g�x�� ������m/B�m�5�:��z�����r�d��T[x��htͥv�OU�^CA�Y���u~�K��+D[���c|R[2��E8��x��	�����"�:�V�;���+�����O��eT�Î���
�gna\�*���:�h�kmR�^l����v&��rԏڵ�ؤ�Rj'���.��>��;G�02���v��S��	{�)�����0��Rđ��?L�Eu����7��xVv�<��9D�����G�����*�� �/W���@]社j�C��-�A�M�%#ʑ%�LҦTO6��^,]V���\T8)��s�-,J�����������C�«�>v"��@�Wy�v)��ً�!0
��@�J��)�(8�
�����zrǃ�����aum���"RWRX���ݱJ��`z�]�>|�8}�;�=|^��&������������Ƚ�#X�M�ÒYX�$�j�j%�0��Hm�ڪcۋ�՘���#�e>������P�U���!���?���ҙ1�X��ta=
�O1CX�b/�����*��	��Ô�DٯQ����i���sO���G��k���� ��ʄ�E�E��$o����q�W::�+�P+�.��%ڋ-?�x��'�������Muuu������O��>�+�?��7ԑD�s@PG���N �EPGPGP'�\u��&����� ���$������������J6���	FAH2�������%IԒ�g��_��Z3A�IL��$���������sHP�\2Q����`����EyS�`{ݶ��ּn_��k��	�.�_s���nX�K[�?ou����d"���%Au�_�z���!ըŇy��_��Z3A�IL����Eu����_��2$�}��.�b���:���LP��Au�aJ/"�#��;T�#��^�[���L����K0���Ô^�?�
�o�'�v���c3�55Й:�N2�'���ŵv�j����N��$��" ��?�.�~�7�*�m�(RGf�8��H�: P_A�IV���k��vS_�~���1J �3̈́�ݒ�M���m���īk��So�����s~��",i��Cۯ�!�h"��7�*�:>P���h�_jf�������g���w��}���9��4/�������Rd]($tL}��#��D�z��^k����j.�Ae�SZh�;�J�����x�Vc����7댽���KP���"�Z�EuL����a��Jg�t :ɤ��.Ü��+pi��lۯT(X�Z�����M�6(�pB`�2���L���C��n��V��v(�8!p�,��a�#O��R(���IF�f8���B��r�zС�^_|���o/A�ҋ(��?���Ae��ui"�Wz�^t(�E��+����HW�D	@�U���%���6\{	u�m�S>���B�թ��Y�D�r�ۋ0\isƵ���Ô^DPGP�w�$��.R��Ơ���*E��]K����Ȧ��e�� k���P�u� E�T��(�pO\�94��m�r�Sq$2�Hep�G�5BP���.�:��B"�K���u� 4��U6�|8o��^(@�ӡ��6��$Թ��aE���z~�YC�,(�%~XQ�����T�v����"u�aJ/"�#��;TR�N]��L�Asib�/��u��z"�-7� c��P���x���11!��27{$1񄠎?<�U��2(�[S�KJA����rQ��@'���Y3�q�ݰ�.��dO���s�&�-<v���XL&Tzn�C���b�P�oC�g��3�	t��b�� ��\��^%�:�%ِ1��q�e��5>_�����k\�&�!k� ��p�KzU����fX�d���3f�u�-�Uu�f�P�(QI�p����&�@O�	ϳY�%�r��h~ܩ#�������0!"��,��]XXӦ�֦{�ҙ5�.BIII��~?�?^�˻��#�q�0c),\�P�ԩS{��W]u�g����sӯ���tIcǎ�9ސ7���+"��7�*�:�P���ta5��!S儂�
�����l�n���p˳����vV���k2�ن��� ��+`��I*����<>��
�5�u�ү���uu���DP�k�k�a� o����Vɋ΋�P��]X���@vI@��=��Tx�K�E�&J�y�M�K�u��x�cK��ʚ��YX$����lt�� M��sf\k����|Ň�8.F�x��hʿ��?R�ʄ%K:Tv��P��xOf�
Y�5Ƨ��*z��=�O��^�W�^Ĵ�*\�@���_)��wH��W�PW������ <��QD5�o�-�������VMwP����♰�,'-qA�b7/uK��V�81��ւ�skjػem><��x~�=�o�x���kG+lh�m���G��:{�5L��N�m���3A�sZ6w(#���䆺���u�mP2���J��=�B�W����o1Gᚗ���g%�<c�$�ݱ�v�Z���+��g����ֵz��j��mɞJ������CE�Sb�"K�ބch�+]�RD���c��)b�%E�jy���)9�,����a�e����=��d�}S�âф�)w����������A?}�|��;���޼9�a������c]�lA�]RB������ͱacD!<�+LPZ�:�oȁ��,��wM�[����q��N��O>|v�Y���ǫ�[V�_L���&��|��S�s�8˔&C�0��F�Sך
�+��(9N�ٸx�ϐP��h�V��`O��hJ�C����xL�2��&q����
�h�-ˍ�ݳ�
~��k���ӏ�Wdݯ!�IPG�:�~%3���>y�s)���#V;���ӧu9Seg޿�~>��?�བྷ`]�O��p�M��u���._R�r����Y����Ɵ��jIĜ9���F�*3�Ƅ���V�4��[��˸L�e��>����>v�te{�؊L�}q���ɓ ������M���7C^,E��V�NWų�b*������t�)R��I&�uYYq�ݰr�T�u���N���'�=���0����<O��G?�x@::�|ߐUqS �g銗���&�2�	�7o��w��}�uoY�[��֮��5Ȁ�*����ll����-���pߞ&-Pp�\ɢ�j٬�|hG+�:%�
_��� Ue� `��њ��s-��=:S�X��:u��&Y��:uk�wD����f�[vB�M��1,��3�� ���~m�nl)���Iz��x�G�?:��w���(1�R���
rJ���.S��>Vt����%�wZ���u����Ȧb;d�/��J�]���������5�>%u�X�ݼ:�=j\��V6�Aes�CwP�q���.��FP�ZHƁ��GO�M��z~.<��$�:���w�@Ӳu��F���hu��ꏶm,�'���� >��o��\������۾��m��xW�˔&��������`(�˙�^�C��sZ`�c4����l�X܏��u�E�Y���5�=��0�!��"��$�~%�#��;T�	�������?V��;��a�@]��lf_��g�#��dC�*՘���g?���;��_�
o�	7�&k�y<� A]���%��
�����nփ�؛V΢b��ݺ� ���^x�ue#[�xAAA]\k��_��M�JOP�`�����W�|7c���Ѿo?�^����gk5�}}w�3f��V�r�o���j�R�B���q�o��=f��3ԱvT(X����g�:�an��HȾ~���>/=� hq�wW�i�uuu: �1�n����w��랉r>;��y��=s�&P�T�V��ן-�;7�0�#wn|�̺���-��=������K!���m��g�k)c3�=�wXnrDO��/�?��:�2�r��B��_�W_���C����Q�?1!,:S׷�_ʠ�Ʀ���TCa0���_	�t�s�q�ݰ
g�(���g��z꽸�Ϗt<��w|��C]{�?b-���̓w2���f����Ϝ���u���9*_���￐XƁ�Ɔ�:��tC��i1��ٞ�X�Qi�um�l���M��?x�i�~/A]�G�ME���z�S׵�0KQa܆N�����őu�8��ت�z��~s/�X�<���� ,�@_mNwj��݇ՆX]@���l1���k1V�J�Zd�D؛��K���y���@{s�uuL�q�][(R��I&�	�\I����y�2��1��Շ��Eՠ.0���`������i,U2�*��6��9Ulׂ7r��|��Πq�.UxX���Wz^c�:���֬�_�~}��{L�h�&�#�#��-$�@݃͑�E3C���[��F�/T�.e�ԭo��Vׇ��4�Jƾ�(�p?s�4s��F�ȝ���e,�Pj�C���Ⱥ���c͙�a��J���W���	B���w_dm�F�i��"uX��L=A�/}�����:�ݗY�r"�F��&���#	�~Ŋ	jէ�z����6�tU�� R�Li��
��e��7Ա&�&yO`�`5Ǚ�_��Sr���8�4��Ð.�}�o���{�aG��OۯIu�#[���`6��9�e˖qw����~�g�%���
uo��n>`�g�8�{A����5{����!���C�%ڪ��ѷ�|Z\O>��iEK��/��n�}�龃���?����`�>f��a�c-ć��̩�j�Ӕ&��X��ؿU�U�ؾL�
��kS�8�n��&u�97�S�n�Uz*i�ף��D����ʾn
��x~���^��ѺM�..�]-O@�F�P�"�����v����U9L������&���%?�O�LM��$[[��ӽƁ:��X�2H؇E��c��?x'{�e�w������SO�8��C���X�-�&�"u�#�����u�O��VL8����N���_�
¸��|��8��fm���{�w�X��{�_��e��5���`i��fy�c�י�7ԉW�U�F�]�S�x�c���KX+iS"\�n�k/=��C���f{�P-�K�/ש�:}��k��j͝�^D�:/��Ev�Pux}�� L�S�Jn`����}�9U�tإ����5V������j/F�Li�D5x�4P�n`��V���&�.�^���c죄�i��J��s�ՋQ�P8s�������?<�%A���%˹����~5ӽ+ni��7�_�u!o+w�R���r��S��:()*���Hg��t�s�q�ݰ
g֪�;/�NK[��9�P�����`�w�jP�3�����Z	|o��8���V�@�ưE&Qͥv���̒��������8�`�����M��ԡj}����âY�����o9c3�	�y&�>c;E�ϗ��/��j��8r��s���[���K��ր��n�]u�UP�����0E���z�~��O�����7�������_���]������{�=�Hԡ�G;�O���8q���Z���}a���kŲ&+��Q,����M�\���p��GրJ��5�e�fߒD�r�`���0˸,��K��y�2�A�b&o����3��{��r��烲��oc��#)d��ˋ���t -$cC����'თ?�g�zv�>�}w2C]��lY�hǶZ��>��X�̖���TY�+�׳�W;�2�?0���A)����o�u���]I�@�xP�9H��
v�B���@��sڜ*�[~^Njo�1���,l�th9Ĭ�>]ge����m��7n��W��,^|�>X��.o!{<�#;}9R�1��-5�mKM����i�����!�6���u(L6������4�S��6�Ε -��ر#��SwIݒ�ܯ�n    IDAT�6y��:�z��ܞ4��bx/�0�������od�.�*]�	���VWP'��B�m��
�8 g��m��5S�PbJM������ٔ"��.񽅄�(�x��9F^�MW�_+��BX�7��;o�Ç��*�za���=�V��V`j���9' ������3C��`�*��~�&T8��ط'>���ٶ���� t�I=A]uYY�kw�X��>i�Uz�2��Q��o��!rw���xᙝRW
��	Y�>BY�.,�3���:���әC�ϚR�Bsj`�)U�2��k����9��a!x��
��2	�T*:��4�c�:�.e�(���
��_	��3�-k������+`Ƕ:)����YNp/0<ԑ;���n�Uz+i�V��7~��}U�b��v���
|��7�A���lha���S�	,{r������:�E�����pkS�Bgz�b���C�))��;�Ca������ʺP�_	a�����<;�'�#($�����u�$�	�>	ۊ��w�������B�=���+���_Wu؊,g��h���6�g�
󶫣a�-<�fx�Ca4���FS`���מTnb+��(�+vS��"}�#�2
T�개��ozqd�hH^�v��h�)��Wo� ��kO�x�3C����G����]U��i��:��|�ٛ��NY[vi-<�Ѕ�e-F��4��#�#�#��+$cB�x-^����aF+�ve�%�E��:����k-9}^Y�&�Ko;:�`�����:�}�_vv���4f�ի�m�~$<`������T*�u��{�������#������A�1�-��}
#�����b��t�C�*2�RĴ�A�4�c��2U�f�`B��ꬽ�~��EG��guu���
h����Fa�T�CA0��_u :ɤ����tǵv�*�Ru��i��{����ڣn���t�:�[�/��:��')��ѫ�Iŋ�~n{������tj\Έ ���N�F*�Ҧ`uu(�HAV�g�~!�Y�O-a�����NgT�%�#�����h!�N]�m뻽O���K�!�Y�냗>�
t?|ѽ-��[i�	c����mV���U�H!G��G��=�'�^n�B�-Sn�!�.��_�L�aF,J�������{� 8N��!+-��^�:�:�:�)���^������x��_^�~;�]�+��ƞ����u�(��<�;Q�½�崵����O{-d�:!��Qg��k�I�4ԡp�9�j�j�_zRc�<سN�ڛ3����������%�#�#��+$cAݝ%�G�G3d�'o|����6D�;���1K��]�+�߬vnU�$�_����,m?]c�)�Hi����^�����]:ϧָuaa�8�Dm���'�Y6�e^ѹ�d*H�������r���"��:�����`z����1������S�¶���L�."u�%%q�ݰV{�*���e�"ޣy�.��!�u�w+nY�߽���"�M��6U��s��┢ij�#��͝�?��ǡ*2��[�v� <b���ՎF����(^��Re��B��3�)�g��T��-�&���8��'K�AA�s��YK��ׂ�u��Wv���y�n����=��}�����P�	�u���nhV�Ȉݞr�x4�.�T�Q~��E���3<愉�X�V+x54ԅ���ۇE7��}�X۳�U�TIڑ��0/��D�L�A�g썕��ea0����.�uuuiF�8��lC�"ޣ�����n�_l�ºv�#|���������b��cm�bP���j�pM�2�������Z���-{�]�]:��#�p���P�����{�����[w-��W�Y��;Ư��uuu�a�d,��Z?��l��WhId	Ϩb���-���	��(�ZK�?���?hU,Ѳu�K�8G��BI�9 �#�#�#�2
T��2������Ov��5/_�!0v=���H"�9 ��HPG���s�3u��&Y���Ý}̡o��������xWkϥL:_���U�A]�NE��	FE�(RvZW����?S/<��=Mٯ�'�[�k<k7��>eٯeW5E�G?z��^��У�޽��q\P�u�:����-uI(A�/�"�#�;-�(�ZHƨS��K��-���v���yǅA8u�T\P��`gĿ]��FP��2����:ԥ�H����?~�b�g/�|;�9uUz�J�@�}�Ǻ�������n�j��a�����o�MP��2����:ԍ�h�fP���AЕ`�$��-$c@���_��.͝\��U���0.2s�Ԧ�c����z�v�wx�ʧЙ��/A�/�"���]�i.���̕1��[5��P��K%�t��8�q�ݰJ��Wuxa�C��)F�0������-ڮP�z=|�H�Ċ�+���͹�D�<A]ߗ�����`�Ա:7�~��Z�g��K��L�b~��U�@T0{r�sp{�P2�1�s^T ?��+A]��DP��K0����Ҍq�����;_wK��M��ෟ�G�C"��uգ���٣H]ߗ�����`�����1���G�K�X�ڦe���t�uxvo��z�wu�!A�/�"�#�#�#�2
T���֪{��)Xi�"E���֔�V|?�t��1K�D�:��w���z�wu�!A�/�"�#�;��ɕ�>gCL�)Y	mMPQVL�: �dROP'x�q�ݰ��P�^�ERr�j�V	�z�=8y�d\���_��L}��#��Bp�JnvA�m.��tB�r�䆼�=R��̡}���}�_�7�����ٛ���YCnP�������|>�8q"̿f�"5�7i�˛9T҄?���Q�Do��P�%�8���5��"쏖�!w�Gjz�u����%MG���^(X聒[\Pnr���h�r�z%{3'�^�C����)^(7�������BC�������@�V�(AZ��M����yi�9/�'�H}k����u��:����>	dZ�l���z+�r�Px����3�� L�Be�Z�mL�Qp@��n)��u��D):�T�0���>`��,�&].�A����fo(��^�:�0���A�H]�
�w��M/��;�?�+E�x��h.��
��b���� �$�&c5ԥ�R��R�B�&��y&��/�����A{m�؛o辰�%��SzQpZ<�}WL=��ؽk�_�Ng��t�+.(�k��f_��|����4�绡�Z���X��"s���Z�o���ؗ�P�aK�ҵ�ܮ$�{�㹠��:11��Y �~�񇦾"*>L5�m��!�ըP�ǔ0衹?��J���x�_�%>hjooG�
��]���p�P�_�E�x��c�CKUb���?�.p:S���&�:��d�����
���]�ŴA�e��B[Mb����q7��.q�v`�Np��B!9�.o�G��DNpX����O����e�<��KP���&�:��d�:#+��ss�E(<C.'�O��L&r��ئ8��{�.�p����{\b���y=���\!A���DPGPGPgl�+���?j�D�K���m_����+;]C]�_=�y/ޓ,-�
[�[�j)0ӫ{�A�w{	���p�$all�ff��l��9Z�l�2��$���3�f�k�vV�B]�5�*�#v��ڞq/X�#{�m��buu���=�XZQh�5�@�0��^�3{���{�H�:�/\��J�PN�PʳN]_�:����PO�:�����_��>�T:~W�h�� �	�CpB��=�фE��^Phoc�>�Ţ�u�_�zAh!�iuX�M�z�j�G����a~U��uh ���P��}�ބ,�\T<f�#�C�:�0��T�*)R'갼o�ӣBVpGI�S�*���u2�'���9.���xп��*^c�^q��f�boT�s�4̊�?Ԫ)�������4�`׽-��s��;{>|�ex�����=wýw���Fe�B0j��$}�Ah!�i�l�&�����<��^޷��۳��{/�[�?�>uܽ�R�R'ju����J��Ze�*�S�Ξ��L��^z�K�2V��k}cC]E�|j��sx�3s��ה*d��|�������-)�����H������g����ȏ�m����c�~���χ~��UM�X� w� �cʠ�Ʀ�*�TCA0D�O�b���9����nXW�p��Z�|�yM���8q�X��觃���n����a�Y5�/ֆS�Ȟ�=m$<bN,3�R�3������.4���%?� �����K��
rA�"�	�C|o����7&�4�X������Z�l�_�c���G3U?���p��rY�k*v�?�2�H��J�PDMoۯT����5oF�l�xz���0�������u}���Ջlѫh�L��k�9�g(�5��Fǁ�S�z&y�l*��kV�v�U����Ä�V�Ʊ��x�C�-�\W�}���Z��a9�}�ٝ ����{�d�78��`	��(�X%�c�V�%��o��lt��a鈐��b�2%���"cW0d��t�S�����Xx�6 ��l���j-d����n��^r(��l�v�;7�|��P.;ؕ.S������޽��!�:v'��=[���]c��P�"u:�A���"a\	�U���K�=��!�ݱ���ޘ`���Dk;H�_�s��/6����:=Ƃ:���jd(���t�?).���V�6�M�vً�1��W�]�������u��`M3[������;;�~%��5XR����g����;����Ӫ���|�V�A%&!���X����j�,i�V)����&y?aMH����:9ի��'3����1F�;E�]�X�`!��3f������5/̖eC�B��$�:qB9T_�Se�+!?7�^%J� t�I=A�=���+8�����/0�|�����=�oeB�u�<�[����S�
���_����o���`���
��@]9��XmY�k��6¿�5qA�!/�����}9�+�nbG�\�/ �9��&���$ꨣD�g���dx��f���!,��P���L�}*�N0��A5y�=��H[��d�5��g�Mr�<�҄�j�Ӓ&\^�q�H��>����w��C;Z��Qa	��,	����ul�ts1ۏ��o���ݳ��i������26x�y!�<1MU�H�`�[�q����Z*�&�y����9�Ps�x��`���80�F΢bm���7�h����cL�uy�C���74��=ul��z6���5�G�﹇i%��'K`�X�{�����>G�ki��`�%�8�B�a����>�e���c͙���eXIZ�a����*0,����7��Q/�%;TR��?����z���%L>`u�K���׻o=ZU�.`KRľ��T�n-x#�Z��L{�A�.�?9# �R�Z�U��}�e,�^�E��[�2_l ��C���0�}C��;T��΁0��VĔwN.dffBFF%J��"Rg����KW���7�I�L>`C�Z]��X*m����v�0�
�Z�F���O� �l�3�BNȊ�n�cgx�dMs��c�L�:uR�����e�����K�d�9��Q���+u�������Aݺ6hua�X&��d�:�0�H]S��H�����=߲���6�@]*{!@�E��k�5l���j�@]k�>�0������+oX2�����/�=��p��ر#����^z�i,�����e�/0��� 7�-��u�e,�Ku���S��M�e�Y�q�%����et�`k��G￪�C���mL㨶RW	�/a��������je�&���k⏰�9�8
o����;��,k�%���VTM�0����N�8���Z�bK�F�2�-j�Ӓ&�Y�R�������<��F�Ӱem>ۼ/���"񝃼)U��n[L�ټ�lX��5t�� Oۯ��@\k7���-I�i�e+ƋY�j_�-i}�y��Lyub��}�O�)U��&od] ֱ&L��z�u�ǍŸ�jd��-��#�q��k�1����+~Xt#�C���-V��쓷�� -���_@$�s@ٯ��;�RI�g���S;p��qU���w�1�#�y��"�������a�+�<���s��E+�@V�f5�h��uN5�hr�B��+6c��6%����>��v� LI�gK��q�~Mv�$��-$�:U���r��ѫ/>��?:y�8l]_�t��J���*����e���{�K�,P�7��
-ͥl�����ئ��,H��
�q�㷥&+v�(��u��K�S�䬽�	
Y����׫/>¼���	�҃�����c{��C{���iv����?z�黙���r&a�G�%K�w�#}�,��@o�a=�o9]A���Ea�����4�h9c���\�����+*g���taa?9�{n\��~�V��ɇ���F�_	��%t��7P�A�S����{bj��;��;6A[S����$�z��`N^\k7��۸?o��hg�	[���?�P��(Q���Ӆ�a;W��Ǭ��,O�����g�^�>�z_�>���:�&�Xc�����Rĥ{��R��s=�� F�05Zɢ�Oe߂EmZ���X���ߞ�U+�3FE�H%��8s@ٯ��&YEu�؟גط`%�[W ��J�7:-��\��t�U6�ݗ��w�G���A;F�~���W�� �����ݧ��QK�-�f]A�7˙���3*Y����M��)!*ζ�oT��#eaa�6%
e�/Bc�<{W59��g��Ǐ���������d�[�EE�yC��DP�n�Uu�څ����Gk��R�9<�����������+�����R���5V	
3�����ׂs�c4�0�9����:�X�G�>�`JX���W_P�*B�U��9��
�T��3��s�@���T1dJ����.�=(N�Ƃ����" ��
��~ŋ
�=[^t2�킔@�u�N�8���������� P�}BV&�q���怠�?�$���=�������iU6���N�櫏�%��Ç���_�G�_)��Og����j�_�s��ަR��7��3��L)b�9U�1������ę�c�N��Ce�[i� ԰P�Ѻ�<�_xWi.�I�?<����_	K�G�:G����G�MJ5�p��Veg�ˮ��!�d�9 ��7�*�:yϬuh��ݲ�BpãB�ֶ(�tV�"eg�#�u�D	��W{��3�8��zFYl�ԥ����SD�Z
 f����P�q��)�J ��Iz�0�r&UĔ�<�feAfF%J� t�I=A��6K\k7,qB9��-����)�v��W�P���W��ކ\;s�]B��b�	Q�*՗SsA�Ux�[��^v�^�:�/\��J����<��)/�7_����nH:���=�����0���-��?_ߡ�0�9����n��T��B-\��pfo۰X�������A��^DPGP�w�$�SuXT?���1(�$�%g<�ݷ�~�
3d�g�+٢_��=;��˃V*]��9��`�<H�N�t
���)����?��괄:�u� �:��*^�]@嬽��R;0޶v(<7�k�Otc>߉����H�֋
�u���lXu{3����	��Ô^DPGP�w��H�r�C�G�UK��+�
�`�R�t�j��ʵ��$�"B����!Qꬽ�ܶ�1�5��L�:�0������1Urk�f���P��@'���ٲlq�ݰ�Ӫ�?o<�.hP�B�������6��e+���=�հP')M��'*KS���ڐ��@/����MT҄?�$����zP>c�?�8����bi!�V!�?k������䁺߅٧Z��W9`�n���N�ImI������콍���?$Mu��&YEP�.�unm�T���de�������^�����r�S�bʆ�:֩�0%�PSs����z���{���e��y|�H�:��d4��dA�6P��J]R���R����f/V�h�T�j<�LP�^CB���(@�_=gΟ��o;b��S7{��R��T�D��\<    IDATm56)���AH2����M���N;��܍�z�y�v����ef�&p���޼�=R�GI�/����N��>u�e�P��^(3��>`�Q/�Rk����o�W��x/9�ëx��q��b�f/F��^��W`/AHҋ�T��w�ԝm�Ö�k`E��%t :ɤ��.7���+tK+��M�P�5� ������POm9�JlR�
3<1��g�x�RY� g�G���e�0X��V],�R�v@�.)p�v7�>u=�M��y1̠MTY��fid/A��^D%M�CI�QG	m�.�0����G�C�vWFS�F'{y�F��:�zs@P���"�:�*�C%A�#�u��� ��)����?���x�	�/E��	FA�ҋ�V��ֻc����`��Mв"Dg��t���ɍk�ո����H����f�:���"����5�(��"jz�~5-7s.�,�:���LP��Au�_�FAAA�琠.�d��W�_�DP���k4����	�K&�:�_�DP���k4����	�K&�:�_�DP���k4����	�K&�:�_�DP���k4����	�K&�:�_�DP���k4����	�K&�:�_�DP���k4����	�K&�:�_�DP���k4����	�K��uY��������P�q@��P����v:�t���y�3�ǭ�Z�D{/�Ap��̮��F��u�_�FAAA]�@]�P�+�P����?�K����j�JnqA�\������߇*�u� �4/,�@E��p��^�Jn>c���x��Pg�@���n�ء��
���'�ӽ``��������5V�v:!p�2
L�%����5�����6�Y��!�[������A��)��Q,��^熆<�3��Re��L'��x5Z�B�}�_���:���q�+mPp�2���N����֦���g����	���p�
�-_��ϟO�9�l,Z��ڄiu��~)�
r=����������΋}�������Tb��3�Է�pP�_�s*Mn7ة<3�z	㗎��M#{����AH�+PG�9����"�à�_�`��?*�A�,/Xt�1�Q������J�؛�P��&A���*���2�噈��bo�� [/��@]��jX۰!�քփ�j�p*s��eߊ�6�`EPG EMP����������S:j���
ӼR�'�Vٜ�����Vѹ��A�ǂ�s
Z��mK�7٧������ѓ�͛������@F͊�h��I�q�O|`w��hdC��-��k�/	�.M�28=�a�=L�HآJ㳠��m���������~u��PZ\xV�yQ?WT��9���o�������x=��+.F|�a�u�����Lnv�y1���AY���}. �#>#
����	���1t�LnN �3^O��s���.���g�~&r���Ě��,G��DۯLP��#����jlgtD��9��[�<��k��_e��[Pg��>q`�`�*����xB]}M%���޳z��G�~�Ž�#>WU^�oUE|��'����wn��̪���{���">WVR��3k:Z#>��wv���f��
����m^�;o�u\;���k:�}�{�E|f�ʶ���]�m������|8�3u��{�6rޟy�����ve�9#����D��r����vi�T���m�6��U����t 8�Ug��n�,rs�������V,AAAAA]�@֔��:��r��v+k�򶳣S#f�)�Ðk���cNt��ô9���D:�fo�l��,,�:�:v'Q�q�͹*"r��#��~�'���\SFG���:�o=�X�����@d��pS�����ӑ���>��ds�g�|_���L���+�6��s�6��-ۣ�k�����rK��<�qg�g������?��ш�vxVw�̾G��L�}e������{����u{i�9��}��ȏ�<�갖)o��U�4����X ��}]������uN�'5��j����Y	�*�������t6��P�s]�����ou����ٽ%�6l�z�nP��{�����#>����}&wJ��2�b~C��ݻ�H�k�;�v���m�[�}���E|fki�τ��V��t�̾G#���l+#���.0�P���n/�����d�:���g�x����D�:g�_���*��}����ߛ3����y5���CPGP���ԝ��:���ס�[��9�	[���{1`���6u�"��	�A�[S:	�v(^���q�D�מ	��=�<�d�q�(�8��j%��̦Z%h�x��m��
�٧������;�|����ߞ�'�����쭰�gt0��4��&u(Rwf(R����;7�¾���_9돾�|?���^x��u��U�V�"�jm�0!P���v(Z�a��g��s��e�os�zNb�
�*���v�f��:�ޔk|(���|�ͩb�)-0589����0���ɔ"N��_�w����-O��
�
�����+�O�����u��	x��=�qe@��JuT�����Hݙy�H���
���G;﬇��xb]'��7^����p�g��[�&Bc�����^x&�~3��u����9���K��Œ"^�1D�3��}Z	�a!dCB�����Uj�k �c�'��3&� o��Cr�
#*����/3Jg��� N�>,�ѣ�����e��Zn!�C���HA�ߟ�ԝ����[��AY�a�
����1�]�ÿ���7ȺgcЮ�l�p�Wv%���^��U�R��72R�G��Ջv�+CB]ɭ.y5�fxO�S��s�9�\ơ�k�������L���9r��l��������������-�V�5yu�Q��áHݙy�H�髪u�G�V59�ӏޔ�N�<	�=�Z�?£KJ�o��=��^k�$�IS����A�s�9��$��b�%N�ui�ԦJ�6hJ��h||��k����
2q�Dh.g������ u��v�1߻��#�#�#���)���sAٯƕ0�DV�{o?��!���V�|o���YCD涣��&N��6�
���F� �#��vت�PP���+��퀌4q�
C<�:ܷ��y/֭����|���wOב#����m�v��ނ��W�~U��P���<P��? �E\���0¦����?�����+�l��Ϩ�,/R�6�l���K���r�P��XP\��M!d�h���~��Te������c�_4�����0��v/|������kO2/켙uqF��͛��e�WTqml-�rV��6D��ƂM�+����t�[����JϚ������~�m��\�U��>S��%�3�j�&�G|�^��s�授�D����Οk����g��[�τn�����e���l���n����g��٫\�9�9ѿCT���9�p����*M"�9:15������.�W������˺P�z�<��o���]lǾBָ�/��*k��v�9E,Ws�����E�g�;W�[�,��{#�}akzy�91_�#���H4��_!��<�k�����?êl��� ���1&,`zs�hU�7c�;Y%�Y���Z/L05�H�j�Ӕ��zx�p��}��l�=u,I���؃k��Qe�]ڄ����*A�㬁�26����j����8��e�_����˼���_�a.+`;3�@�y6�h��zn��/,㨐�,��$���k���l���q�LL�4)�u�e�qY�hh��m�9���?:��O�������i��؃*��ض�1��9XxYm�p�����l[�X��0P����<@xF��fz�������Ůb��ŭR-.,^�2��r�g����ӓV�G��76 �hh���	%L>`M����\��(�.d뚁S�x���7�������`$�:+N�Z�U��y���4�Y�$	�.l'�2��\w̗��so���"�`�Scƌ���fr��i���L.f�;����?x�i,U6v�����lM)B���{��c&��8uil�:���Ok1Vq���I�B��"u�5�N�<��C����0�#��#�#���H4����ar�V����4��Lv����G�R�۵���y�X�R�� P'AN5㙺�>M�7��֋
��x��ǃ�h����^�q�ű�HPGPG���րA���R�3uX�T���!��2�A)���q�������O����&���^n,Ɖ3���[���TqB�U��f�*i����#��Q�;����&�~��W�ΊDs@k �5�R����g������4��E��A�"��{O,��5y�T�:�����Q����He�Li���83
XS�sf�[T�u����ЩS�`�� �8Jg�|A��j��nĈ15j�(�i�ȑ1��sut������ր�@C6[��=���;"%a��C�.�N](�-��2K��DMް��cmU��@u�
�w3'K�.���/5ƈ�3��T�D"�q�:J�s3W����\�/��gc� <c�:A����^�9Z ���)��ض���`��Z�� ������-8z䰪���Wg�G�Q�:J`�/��`�'c��[|��µ|��/�E����y@�@VJf5���R�^Y�-M%lQ:�e�~�L`�w����=@'N�-�
�@���8z�~�hh�Ps��c�G�>y�j�����RV-k�ߋ
�bm�i���`�':������Ul��X`��6�@]�@Zk�&�`�i���4�z%�3���Ll��P�e,wQe���KE}��˪<D{����!!v�+��� �Z�Z���^��V6�����U���GX���)�ѓ���̵qq��=�w&\��7,i�f��[r��XP�������{��(��������/t�`�/J�R�~~Xr@rM����}E����f�/���\�/��Z��_�~/�OX����\�?z����o�2��5fY��RnG��\�����%�:��H���{��:�$�E;q���9U�X�'Ͽ�3�[��=c�P_r3;XI_n�,�/(�g"�l�>x�%Y���G�=��3��)9TZ�h��5Pt-�l�>��o��k�>��fY�ĭWKe�7��y��҆�r"
��9�0r����M��5�ZQd����pС���������T�mJ΋:�~B�)E���x6䱓zX�7�+e�U��c��������������
��*_����!���5@k@��MEr���|t������ѧ�	wl(�폂�U��������:Ӳ�:L���O�,K�)*�����_(�{#�ɵ7wn���
�P�4yѺΓ]�tB��i�8�G���2
[�	�{'{?-X�a�-2�9T^�MW�/Wf��F;���
o��W
�cF�����R�W_|D̅���ͧ�)9TZ�h��5�7W��QX��R����z~��)���Ç������?wnd�`�U͘�:H��uߔ�����V'&^�v]�ݟ5��0�m�o�o�����R���{4��% 5,����N���Ǯ�̢j���l����\���pH4�h��nd�Q�{�ɭUi"4�)����zv_�P�H�3�FM�p�V�^~W�G
�^�߶hj̷K��u�Lə��5з�@֠p�e�M��D��2b=�{�O��ָ�{���P���{B�mC:F�+6K9s�g/���3����hh����}\�V?��D�m�o�b���-��Ul�0P����϶$���P�BKef��������șP��5�P�Ѱj���o�U:���M�c_�����*5d�c����91��{�Q��U����^����_j��FP���K�9�5@k !P��h�u�>�o������AX}á���,� �k�Ca�O��	�>�Z/��������KPG΄��� ���:	t�|�.d��y�]X֡��9&N���=[YDR�P'�Ny�&]��	��cm8�V�7���A�.��� ��DB���Pi�����®Mr#v5+�5�l1��$~щ��b;��ks(��^�~���-���{	�șP��5�|P'�]ڙ�n��?����΋�)SCa{�eo�]�$LCA�>B��ɐ�u�:O����~�����f�=ˆ����Ds@k�� ��1�5�c����c�R��=s܉��p�������ԝ���.i��^H���u~���f8����ܟ���	�Z�u�(�0ͫ��gWa�t�K��%��&B�J�T�VM�+��6%K�,ԅ��z��Tʛ�Ơ
y�v��������Pr+�+o[��/�p6{	���pI4�h�����L�I�[���#�搿�-�[��0��r�S��(̮�mݬ����Pwv±��X?�_�"n���ŵVڤ"��6���X�! X�FWJ�u�O*��U�h��^�d/�VQ�+����	�Z}{�B]g�gб� �g;���v�abE�Mں���"J�(Y������%_�锢�x.=l/��� 
V�����L/X/L��}�H��A�.��� �]B	�2u:�� �:r&�h��5@P��ך	��Ob2�����Ds@k�� Ahֱ(R��/�"�#gB@Ak��@�^���k�u�'1DP���K�9�5@k����?4�X����`��g�AMu�,�R�б���d�U��I4��cP����5���d�ޠ.���F�
o�L�X�<U���'���H4ɲ���Z3A�IL���v8$�Zu�}�Y��W|	FAA9T�*Z}{P����5���dAAo�C�9�5@P���u.����K0���ȡT���k�"u�}�����$&���x;���:޾ЬsQ�N_���c��5.?B��A(--����E����
ڋe��5>���+"G�Ck�� E�t��:R��:K�c}����.�8�����6h��BK�V١���e.Ȟ��?�/@����~ȟ�r��E{�:${sf{�>B0$���s
\p�p��'��O�s��9+��'_x9tr�h���Dp��Ap��3�P����~�5W�`E�j<(��ٳ�`f\���_�,�@E�B9vh*���m�X`��JnvA�L/X����Iu��~([�&���ʬ�,���L�R���$Hk��g/>X׻�6\0�����?�����0h� HOOO:�=�M�&ݤI����#��a��ɡ��5��,i"x/�A��m���QC�.�`��G��^�dTX\�V#��P����z�v����{�蔜�����-Np���׃�r�	��m��BE������s�9��������x	���8u44�x@0�+E���Gm�V(�ͥ�ݳ43�А����6(�եI��pP�[�5.�z0�0\�9H�I���	�7c��{�C�{�Я_?H�5
��?���ԑ3'��5������V��z�1>�5���*�Y$)��>�ܰ'�p��\Ph/��'��R�tF@�P���q��Dh����������H9u;Z��:���]�"j��Gx,�y1?���=Q������.�!�%�>v"&��pc�A�TQJ~H����s�zu�����W\ѧ5bĈ����ɩ�S�5@k@s�������Z!p�7������6Dp�S�}�	vk����BV^�N؂�$@����(�.�첈�о�1c�D��"u44����e�/�z��Y!+��K\`�:T�P����ٳ�}�0b��:+��`��jz~��E>Huu���0B��:)`���C9��mWv��:���{�;Ot`���`[��.,�:�:��Ds@k AP�&B�áT���d�J���z��;�۷�.�j�����o	V��џ��v�䌽uu�P	�h$�aQ]����Z�l��<)Z�֟��6Y��t	uX+����FSC�C�&UsA�G
ҡP޶ESc�.%����v8$�Z�Cvf³]�}Omi�    IDAT4Չv)������z����0>�Yt�&lͥ��KX񛠎��*A������@}�c�@�]-�|/,0p�ۦ�^Ě�;��JՊ&!d�����v��}�u��;k�x��"����O�<R��۰�C�i���S4���vص��ys/|���p��a8~�(�v�g���ൗ���T*���������W�~���H4ɰ�����UMx�����[���}G���G���>�/��wn*Ut�k�U"��X�N�X��P���,�i�����C}�H�1\������z��V�=�JmLŉuu�S�z+#�L��۔&�u,��S���^�9�[�r�Ux�K�EU�?��\�~�����~{��{�/��QI�N�Ds@k@�5 �-��"���O=�	~��`\�賏��6��G��*�F���\*�ސU��n&|b�'Z����7L��g�
�i��+dϭr�z�	u��!7r&N��6�������x�t�`߿g�%��{Vڤ�o%��3Q^�nM�>x�%`�N�:��Gv�N�P��J�:�ԑ#'��5��(�6O�oX���>y���<y�zl���³���Ȏz'yO�S�C��o���O���&�=Vڤ��ᠮ<�)���}GM��YcK�/��uB�D+�v-��	�W_�J��_�-ka/�!�����\	�h��5P�g���m~�؏�k�����o�2�[�s��Hu��Y҄����%��,��uZ������%�e���b-5�
�i3%�C ,��=bWew������=����/���'�`�wH���J�q`�(JrL�qji�
L(�>fRr��M�n��n�	/^3��	7,��G	^Q�1��C{=�?Z�h�/>{WotZ:J���-���u��9�kǹ��N��𕑖-�i2Pr��XP�ľYnv�)U�Tc��C��b�=o�2���Hݬ��޵ԺN�8[��-�Z��ң�W�~��vn��-Z$i�ԩ��d�7o�����ɓ��A�X��$Y��@��UpsE\�:�{�of�u��7���06������%]~�彮Q�˭��(�Ͼ���w��0�bcG����e6�P���,�����o�Fx�ú{,�ǄCAf�0F�i�;ۀ��Rc�x�.�*�!�/�=N^1D�'�r�U+��@���w_d^����	w:uƅ��9n�ܜ)i��7�ߜݣ�yP0�V���H��Ü0a�.�.�z�4�p˵�{��BGߌ�&����*�Í���uʖ�1����]!jʔ)�~��#��9}Ҍ�s��ɽ��e˖�8�8PW�)0���-�҂�כ�>�����}j��A�`�{���?�����R��}��^�0�p+�Ÿ�,'�RDA�qf�����9�V6{1M\�'6�d�uT�8����u�F͊����Z�����C����y�Z7����j��ٽ�Cm����_�>���V�&�O>�7'M�ԧ��!�-����-���cǎHg�Y�!N�w����F�RXR�%j�m�on�}�P7P�Z �L�����TqPc�F�M�R�r�����>��z��ML���'����];u�A���bL�%qC��7ܢ���R��4 '�5�록mL�(X$/��z��=�{\�]��eJLeM���z��:�Iv��i2���,��e9�
ӢY����o4y��h1�8�^��&K�3�[��"u�;�Y���;Rw�UW���"��7E괇������eef��7/e���|�͚@���nTM�-���?:r�WM��+/<�4���{3�m5c4-s���ڬ��C��I��-q��
K�^-��Oi1����,��-�d�R���;訪t����}o���}�׽���w}M@T�IA�AQ�T��P��9���0¤�$*C�L2�0*�$B9t7������V�J��ڧΩ}N���_m�����w���o���)|/��1�}|���(��t2uօ���=4T��ۗ��7Y(�e>Vd�M���>� �hK����ml\PW��W#�CێAC��������},h��ׯ�
KV�:�?��:�Q�w����J�=2wM<[�����{���{�r�E����G�SS���5�^��*�{�sjy�� ��Z�Q��㹗yƬ�hH�:�B]�6=���޽{��N�"긂x_23&�m��.�{p��<�o��N|';�.U����G��e���R[�A��Qv��F�F^�y�˸��H�5c��UF�kN�i.�JӘ��̗����5C^"Z�s%
2u�է_u�:@]de�h3�Q��w��,����w�A���j�UF�F~_ǗzO7����-�Υ�u}f���R0���}��
-PG���=t8���#;��c�k� u��P�(2u�ԙ	���W�5uW��ҐxT�o��k꒚q�����;�z�Fƭ=��t�QCց:�ݠ�=�lx��V�ާ�=oi��C���4-�o���c�y��nX�u�g{0��L�V����9��W�@i�8�xt��aC�����s�G� m�'xK�e=�yC�KΟu�&��%9|ܓ��B�_'$���d�:�Y��}&ߕ5�wZ4�	murxϹ%g׻є.-z幏1�Q������_���:@�٠�D���л}w�k�`&�����|;N� X�����]��:y�2PW8��؎��ͺ�=�n��������i;Q����{�D�'�Q�;�����
�:d��2u�2u悺�6����o������
�xd�Wۉt�*��̛��R�?�'����r�1/���e���u��с�,T��%���u��[�-�
�u}s��՝�Z�*�~wof�n��}��7lIߋ<wR���P���� 2u�m�L��lPWԧ�;����W#@�=Mb���B�'�_f�4ΖA�M&�
R�w��j�r�&A�`�7�@�-�� om���lW(�'5u �~���7>����#5[B~�nܸ�6�+����,!�ꑩC�N�� SgN!Sg.���];�t�������?��֭���ݔm���+��<ǒIq�Px#���$��7�)<l.�Ӑ%Q����7lqre�8o��m��q6�4(�9l��E��Οag�N�	�*����^�Ⱦ���0f�P�$�`�p�:�CiJ:��M�~t�n놅�④c����H�7����~���d-'H$�!Ϧ��7���zP�eJRU	��`���[96�{J�Mi�|w�f��=6UͶ��T��w��M�խ�?��3����W����hNq*�;��U�L]���ժ�4`���#�P�C�ᐂ8��v@�a㡮�w���@���ƽ4��_�
�ݮ�(Ҿ��#�d���M�ej��0�I��	��b�i�]�)|A<�]����TPG���Yj�sSi����۔ytX.�qݹl)V��̵8���'-ӽ�F�PʣI��<zk�xv�����Lt����J�Z�k̐�2	����N֤I�hтu��Y8�!S�k�(��N ꌇ:RI��xDS��O7
sׯ�����^)�_G�Q��hT�
�Q����4��4�|0�;[�<���`aL�o�ych��I�U�Jl��Y���oe��Ӿ��:�C�����CL�y��p�e�Y'���$�)Ǐ��t�v�z΂Kl�m�M]9:j�����Yծ7��S5�S�9���.2��3�������W�j̀zmq�-��=���`�[������h�D��|ӯ��ԙo���ݕ�Z����r���A��'��xt���j��m��s�!����B��$���l]���秪��䮙�f~|�72?��ф�t�ӣ�~׬�頎D��jh#��=��tu5�ƿ�.��y��2ZY�(G��ԑ���ԩY���C�.`��+2ua���f�lR����q��/M�����T@��	�6��.�n���s�D�á���U�]��ݷ@)fꯕ���{�m�<j׮�pp�� u=|0�>�Km�b�����h��D ��qi��[����kJ�#��yZRox�ܣϴk]��N^�}���b���7V���o�=h���u��P����u4�+�B���[�ƦU|W�r{���3G�Y�r�@i� �S��<��3¡<*h��N�M�F*��u�]��P��E/Ե��}�k�l/��uZKn�&���F�_ʊ��g�/��҂,ab)��i�q#�;eД.�����/��/������e%�kٲe�P׶m[���3�z�y�6`>���ںO�>lܐ��%ML�Q�� �P�.h�sd8�u�8���Lv�Y��P����	�MI�]���aj�S��6��C5ix���X"!��o#���%�yLAUv}k!v瀺��~�M1�TP7tЋ��.������o�@�Pg�ۃ�̇�t
�Ɣ�Y�~���	����s=��E���l�]ؕN��̇C��Σ�ga_sFk�B5�V�w����w��e>�`�u��;6���֩S'ᙸH/i��'��������/̊x��	�N�S�34Bϵ���nJ�tà.-5Mw�{��#�T��W��!a_�N����r�'Y����RYz���k�#`�I�00ms6jSD���1�ٕ3Օ����jPG��y���`���u��E8�� u�:@݈g��#ذ��!R�gTA�ȰC���E�<�xDE��������ֶ�kWo����RPGJj���AM���9RX~_���96�����Ɗ9Z�<�Zt<qLX�e��z�,yh����JLy1?�r�����	2u�g�>�M��F�+S���'k?��,?O��Lj�H��2j�l�8;�y"S��aZ������AY��cS���yϖ�:���[��24�H�-�-{Kِ�&�k��PgeY}�u�ϳ�{N�_���F�?����A��<xp�����t��k��=�\�O<�D�P71w*��g��e)O9U���fr�Q��;�u���y��i��j�3s��9'�h��5��l�p�`��:�+�Nj�[tN;�-�fg��%�r���jY��(���g���mpZ�IiOJ�&4�8��R�y}�l����BѶ������Z��:@����s@]m��[f�����6LHNg��Y��e����X� �z�<oi�Nˢ�F���P�-*�GG��e��?���5c���ؘa,���9;�L3��T4�s��R��Ɏ:��HWw�?�T���H�:@*�
>�>�u>��\��G��7U�Gt2��٦��Nu�U@����%S�/KY<���i>��3詿�g��7"
� �l �ԉ8l 0/�A�)l �3�C��DB�}���]WF�҂�H��w���w���� �Lm&���
	u�uy��s�=�[n�*M⽃.մi�z@��?���� ::| > �3A|��H�:<+H4��8:��7��MTC���GֵkW�bgcπ�`�@�� �_��Z�N��Af��nݺ�;�����J����[ٓO>��P'> B�A�� �N|����1$��'e�t��N�O��OQu����g�]�:��"� u�c�P'ވ� �P׿� �񁎬��Z�n�B���#�Ϩ+��
�3k?[��jيu����D{,Ix �`�@d� �N|����1$��*��86y�dn�7|Ԥ���IRi�8����5}�X���VA�| > �gm�:��� u������d�/	Ň�?+P�p � > �m&���
��PU����d���Z�N��A)��Y��E�P֣�4�O�7���պ���~d����s����^,��l �Hl�#<�@JH6��L]b3����Yj+�zذ�nL	��<d8����>Oۦ���?w�I�>7�E���s����2N��!� > ����f
K�Kf�����u��P޸��+6�Fԥ��b�O8�8)�M�Nes&�Y���z�5�Φd��Q�g0��Y��vM��[f9=2ٸ��4V:����z���x��=T��?6��<>@ �������YIN*�;�~<�W��f�����46j��eu�RV���V.���Ɋ2XIn*�;9@G��dG98�e>��o7>�Z��@�HS��T����D�81]5�hGiL	M�C��Lce�;oJ
+NJW_(���*@��g �����J����dS�TM��T:9EA�Y��o^'�������l�D���˰��$���w�9��g���2|���<u�x��
�9Ԭ����_�Ι���+@��g �������)�`s�i�TW�|$Ӕ07r�#�lX�FM�4f-u�a�9R_��դ�tu�hg"QqF��_B�hrF:Kme��#@��g �����J�ml<����.��W��-��k\畤�S���0��.^aE�������������4tv��J��9,�"n9:4����
5}.e����{��s����������Z�4�Ō��"5�N�3���xDk�h�4\��]lgY�fE�%7W�TY�<v(�	a޵�|������C�K	����@���nY]��XDY��gaN�{\lFA��[V��.��x�K�Gf��~lL���d�==?Ml��vzz��@�� ��9���N�i���K���q�YN�����;"����<���R�F;T�b~������g(!� > ������"sģ�Ì���{d���)ZzyP���aD����8s(���JL�O=�����u�Е�+Q9���L3�:=��|YDA'm�z*I1�����&�N�7!� > �X�h�Sx���y�R���1�X��_Y͝bg��]�u·�¶�WT+N�S(]����qvu\� ��� |�x�Z���N �tp0�x��-Sx������n\4��4�t�Ҡ%)l�x;�9*U-Q���G���d��J��Js�ْ2��x���R����Vv���� | �}�JyP��#n̟��^���V,.d��8u�Gzu씸�+�8{�]=�߱aZŻ#�tPGǎ�b �rM��x8���f�:)N)�b�<[�<�~o����ꄤt�����*NLǜ���%�d�o�j�t����5�ݾ��[�чG��M����B�/�=�@�| > 0�
��h��v���}�>�~��G�xt��W��Ӈؖ��U���Lz�3YC��+�i�+	�)o���i�R�<3�Uֶ��&�i?�Se��|�e悺x��M���?����&�R�w��e@���'�)=S[��&��5����P��Ժ�� �f�zv��,����W��5�w��l�	�> ��,�֣7�v�����~�T<����ƵsB��G���I���NNa�}�÷����4 f�o������b����΅R{�g�����*Hk�0�q��X�����[���[�8yx^o�u-M��Hp(N�ꜥ����~Ĵ������w���RXrs��=�B�| >`����i�ϕ��5D�*Ο�Vc�C7���i���T��Z�R��{�@��
�)!>[)�q��*s�w�=�u��:5M�!�����w)>���{Kh�z@���Z�tln�жXk���/�����Ο=�)��o��r6����|@K	1Z/w��/C�G'��S׃�~7��J��l!�K�����8��ޠYļ��kZ`�6�X
�(�V��Y�)���I��CE�:~�5������Д1��-���>�|��ю�l�v*z�1�"������򁔻e�X.�x�hv��]���r5w<�`�S[���7w������f�m��B��c���o˰�i�FM��l�r��(5Ud��+h
Vk
�����w�^�ƍl͊���w96���b} �;�����ͺ�#�T��Ց\�_:!�)I=6d�,~��_�Hj!ϦYF���-u�𑗚������h��k���Ag>�����v-��Pw���>���cU|��������V��~�1�M��3��G��#:ߜ�F�2�m�>�5��Ŀ(�{:�[������u�2ҹ�b��(	z�gB���K�y���3����ߝ[^c���#k�@�| > 0�L��֗�\�{4�lݫ�\\���Cۺ���|���<#�i�w)Sy�ٹ:gZ�f���\V���J��    IDAT_r���}ޚ����(�K.y��ܙ�̈�gǪ��r�`� | >`���<q��ѶnX�ut�&w�6oJ��Aʸ?���&���'o��S�MJ���N�@/����:kĽ��u~�s���kΙ��T_�wC^�S�Σ��v�� � > ���T/�'�N�k׾7$�y�/�0�?�@��xג'4�����z.�k����:"g��7%),!N�jĽfww�12������|��?�d�Kt��ɰ���`� | >`.��
xb�+s��Q���{�ӡx�k�����Ʀ2)Ny��������^h&�P���K��H���q�r���FCN/�N���ߌhT"���(k"~�`� |@/Hi�9t��Q���#|P�a戎���:����1�7��8.�]��P�%s�x�RcĽf?�8�s��Aˋ�;�|��w��D�{��#3	��� |��ǃ�Ā��2ԒXF����9 '�?�ҹ�<�QZL�D�5F�F~?�7<�2f����w�f���_��F����<�����h�"���z,Xc��i1:���� |��>�[�ߨ5޴��r^�0bI�-�N��܆6)�_���>F��M����������)�gw���ۍ2r�#,[�	��hו��Tl ����3����N�7$�Y9),%�x�*J�L&5ͼMOް��/�V���i�ݯ�	|�:M�ŋr���i�ϵ�6ap=����䌓���z��_����-���9O�v����s���4������=}����g�{j]M��{Rҙ���Ύ��x��|0�:PG�7�����z�cbW�Qϧ�lD�g��ż�E;U�l�U�����%| �`� | >��=�w�����vI�x�{�
�{�͆��CKyO�����֮o_�����!5�~��T�:3�2P�ގoG
�$7��n�w�zT���up����C4�Di��(��ұj�m=�W_�M=�و�� � > �X�(���ߘ�ۆ��}v�-��7I�Bh���'g���xye�G�ٛ�{f��|0R�%[���4PGe>�xM':Hq��n��;�%�ǆ�q�m������+C~�~��:������ȁ`� | >`�ļ�I5�և�~��*{�Ց��=j��#+���W��=�!V.e3fʽ��T�����qX�r�YA�SVdܚ����c?���+x��=rt�p{�o-�{��\;�]��������_6�������fn<:vh�v���*[��dMߛ�6��@T��{KRXn/u��<4���ެ-%yx�$��[��uT�wk�G4?��<��UwO�.���L��}�ь�T5��S�[������tF���iW��	{s�xM�7s�]=�C����� |@ȸ�	�G��-W<���.��2t��������,i^����=R|V� p�[\v��G2ݳ��gIT�#�~�
�HTM�c�gW7\$5��Hqr�->�v{S�?{�r��fR�����UMS�Z���C�]�T�N�=Pe�c���k?4\������v���L��ߞ���@���"�x��ֲE��ı�F���+��]�,e�ghK��\���5�--歙�R).�Hh&o��e�lk"���|��υ���}�-6��x ����t�S��ϒ���۸4g�<�7���E�*�(ݝ��n��C�$'5$㒨��^Y���\ܧi���MS������U��Ӈ�����տ������yG��5�6�������CV��q��T>�|w#;u|���Av��.V��M����>�D5mC�%�(�̐�g�$�z�T�@�7ndo�q�������G�<��O��:�6C5���|Dߵe��St���1d�H ��@4��xI���*IQ�S��R:3�7�]����v�h�����Qg����VQ� ��� | <>��\�>q!\�����M�Gִ�,9�����:ϢM޺qF��� ̈���Ѵ��>z��:�m�!� > �X�hA(k΍���T�x�1��օ:�\�����4-�2-ԑr�t���D�T0��)�{�����q6�����-�<��cS�.�U�&Nt?˼*�wk�SC�`�xCS�B������9��sl ��"�F���t�]��
GǼ$��s��Yjk�	$�C]�/A���t��X�N]Q�o��9;"C'z0�`� |�>P���3�Ѕ�H����\�2�3tT#�>X�Hr�Lu�p8<=?5$b���ds&���TP9��N� 
�����| �LM�j��i9i�~����&V��]��)WKB��ĉi�ڋ+�U2��t�p����JqD��J�m�`� | >`m���Y��x4-E�)�(�6*m֤���]I�zD�^�o-u����;���$7�T��(��өγ����i�N'���h؝lD���S#|4���bW��=�
I��9!ݟ�y>��(n'6�����7�}�4�D�L�ŷ	,�q������������c�f2+��P��uq��Tu�S�J�z��h��p�N���5�.��;���V#Xbb"KJJ�Q�>}��?�z������!�_���,���������(H�SV����)�@S�TVĬ>��Bf#;tI&�+�S"�u?���P�_��hg��+�X��J����(�,�i�V�²:e�ӥ<��#Q�\�o��_����cmڴ�'@�������w<r=���l���8�Ѵ�����!ow�N�k�zF=Ж��B=�P�Uy�����Jm%�F��)U�� &$����3��,��S�""o��O]j����`ϻ�y��7�"�ԉl �h���J3@��KɖbO<zޡn@�e���c	񊺱P�Ɋ�q��PT�H��_�EKKŨ��,�qPY��:�� �����5}@ԉ�>�� > ��l�:8A$��E�R��g��۲^�u�H�k�������=6����.������o&��smF���l�����5�Y���ζE>׎�;�������עn��艉>�g?<�������ѦH��@�|@�2uxqL�� �"G-f�U��QJ�܀��1���ʊ�~����|�_3cU����x�ϿY]�z�k����s�ا�ASݾ6�S���s��-���%K|�__����7.^�s����^_�c���v����
� uxqL���j��׬��!ݟ�q<���p��i@������P+_Ã���<s�0�@�Խ�*1�&�y>K�Ň���P�q�>|@�<�����x�x�u���:@�h�`�h�),P�Ȣ;
Y���E� u�:�>���RX����;[��]tg!�� P9��D� D�H�:�I�r�-N���NC��.r�ԉ�A6�6��u�6�O��bI�UN��<d> �"G�:@�h�`�h�)�P�i�1�����^R��h#@��.r�ԉ�A6�6�DA�w��凤X����mH� u�ダ:@�h�`�h��P�i�q��Jq�[�r]�a 16 �5n�Ҕ%lÂm�׎�+����}�i�����{{�ϵ��;����}���c��4zO�+}��Ѫ��=w�ϵ�W�x����u˫;^��|�ϵgN|��}�q����m�����|���V����<�s}��*����VM,ǘ��> �	�<M�KΟmqr�-V�R�� @�يo�����n6��ǫ?�X�x> ��<�޴��m�r�'_m((<6@�PX����:İh�ᒙ����(��-V~A�SN�6�C��� ���%vKV���;f�=�cd���_�Cd- ���%fKV�:�x��F�T��$ڈ�.�> �	��l �C���8-Y�<Mj�y�-N�.�)߉6&���ԉ (�l �C|���,Y�<-!��_�YC&ܩ u���:� Y��:�c;� 괴����v��b�p"�H���D y6 ԉ�!P�Ǧ
[�| �d�
P� P�� P'~l�@�^ǐY���D y6 ԉ�!P�w�$�형b��`�|� u�:�  E� u��vH��lM�X�1k�S�����e��D y6 ԉ�!Pgt����y�2�2�/�P' �ȳ�N��)��p5{S�?�1d�8�8��!Hi��c�L�!� PPB�V"�N�^;fmq��q�,2u�:@�1r| �: `� ����2n������p�Q�~m�F(>, k� P'~l���� P�@c)N�����L���l �$!6+�:�&�ɓ�8�:@  im@�-�\��kP��$�E�0�ڸ�0�* k� P'~l���� P���*ሀ:o���� ��:@b���~�!SW���( ���d� ����_uf�_��_�Cd- �ď��ݐ�������!� PH$*����? S�L�ІL�����$L�"S'�	u|6��+����W�c5����:@�p'�� ) U��?�Bַ��L2u��P��� u��_��6� u�:3��Pv�}��6m����?�z����{�v���0��x�6��+ ��W�c5����:@���/�C�N\��e?X���,�F�:@�P'z��S� P�3� u�: ��_ŏŐ5m a�ӯ��P�g#d� = _d�D�ՐbJ �bbb�\��??���?�՘^�%g�Q,��zW�p�ԅf#@�P�=V�Y���c�3LJ��7��bbb�n��h$���$����D�Pt� ǄE�V�]+���aR�}���PgaM]�6B�N�@
Y��:�c;���WԙGn�=����G�Q���P' k� Pg=%ޞ��>7M�6,yG�Ϲ�$d���f�W�Ѥ����	F�ۦ�|W�����KϿ��������.y!�_Fˑ��f����:��d- ꬧���XEE�&<xP�Ϲ�$@]�C�ѣG5�(튄���N�;Y��:덝�:wP����,.d��Cd- �ď[�:�!����L0`��z(zl �?n�܀�p5L�b��JB�N<$@ֲ�N���s� u�;�ԉ� u�<]6 ԉ� un@�P'z`1���	��l �?n�܀:@���.���wU�pU�l>��o6 ԉ� uE�(�5u�B]�㓙ڥ��� u 
@�9} �:�	%M܀:l��P��!� P'� un!c2u���,.��� d��=�ܦxu�:@�	,@����`��z���P���Ɲ ӯ�+@�� E� u��-@���F��:d�,.L����Z6 ԉ� u�:�41�	��?X��y(�l �?n�܆�62u��!Sgq!S' k� P'~�Թu(>l�L]�c�k��.?�:u�:��^ ��C����Y����C�Nx0�`@�x@Թ�0���W@�Ņ�W�
`�:����m��P�ԙ`�ԉ���_�'ԩs�P��q'�����
P'>�C�e@��qP�6ķ��C��:�ӯ�!�� u��-@�P���;2u�+@�� E� u�ǭh��˗.���`���a{w�c�;ְw�6���������!S�L݆Y����]W�m�N~"|ԉ�l �?FE�]fGU�u�J����lz�_-����X:��߻�]��1����v�WG������jw۷�mv�z;q� �|�R�d��� ������w���rM���	��p��a����A.���SXͻ�t�d��:�5��5�Oeg���s�������*�+@�\��M�fiRJ�\@�	;��� h�| P]Z1v���H��
�`f7�yk�2v�Rh	@��Pw�H[�0����p�PX�u37��� S�` 2���:�IP�g�ڐ`�[�g�4sg�{!&&fD��}���=��lۦe�l�]�%�߻kmDBݼ��l����
ӯ�%X� u�A+R���{�l����~t�P6��l`�n���]�K��d9��ټ���r�ꈇ�/bbbX�TZZ�C�̶��X7j���p����_�Cd- �ăV$@eԖ-*������S=gmڴ��{H>�v�tv����	P�3��v� md�l��O�gtc����l����/6�o���g�7@��P'>�C�e@��q+��v�����Ӌm��N�G�۷c�r��ݎ-+4��+�d���?�ꏿ���111�Vdf�>:�-����M�2�ޭS��ۻ��l�~�����ny��N����腺��G��~4�&�'||�u֕��ٔ�i�j3v�>��$���e4�������J^�L�۳s��<�h����Fn��;�)[�A;h�pJ@��P'>�C�uG�gfmS�	_"AFAݛ�&ԋեӒX��m��:��iX�c�e',�NG��B�����]]�������f─:��N|�����:��V$@��E��buI��t$9c�߸���{B�N?��7�JӮ<�m۶l֤�z���Q�8%�N������N��	P����b5M�>�@{��?��%?��4M�M u:A�Ᏼ�!��>a�z���\��ԉp u�<]6 ԉ�"�6W,����D��k�G��7Y��HM��38S7QC�n��������^�.�T�S�'g>3|-
�~8!���> �Z� u����fNJ`]:?�h��������g�����{ԅaM]�ԭ_=��P��8!���> ���v�Z�����m����.��K��A��������˳z��Ӛ�	P�#��	�ʙ�������z�zGDB�W��������c%�Y/��F�(a�V�/�C u��Ň�Cd- ������l�\�V Թ٩�4x���#Xjb6tHO���'Y��������=4��N�:u}����SGӰOt4 �=�T�@G��Қ�H��C��g���YA�),�l�uae�knܸ��Ll�ޖ�Q��א�8!���PWj[��}�K��.�w��<<�Q�yr:��&�
un��ռ�U-A���M���{��|�ā��>0�GC�H�i��R����Ύ�k�3����M�R��l,�Q��W����9^g?��s��8!���P���_��f�AA��5���R�*`�Pg�s�����آ9�0G��n߼,$�#�t?����ٰDb'QAc#1�P�Z�[~�M]�;w���q|��,���z�\y��w��N6�"�}���l�S�j������� p�s�����6@�u���v��gN�5�O��+��.��@�PG�M�yk�����jw��N.�����Z��-~z6�<w�����\K�7��J�_Ȯ~���7��}��,�hYT����f��>@���	�V�:RY�r6��zcZcP�0}�z�������ZP��E'Of��%�s��Es��������!g��3�n���_��ƴ�q���p8_���Uכ>�m]���um��F�d辽r��u{^�����G.��P'>pB��U�neQy�1�1���t�ֻ�	un/�=}�;RŪ���.�:r����������Pg ԑ._����d�V��E�ϷS�;:
�~8.PGS{֧�f�x5��Ip��2�x��޿N��O{��o�:���uʏ�3�,�y~����h�:�C�;��uޢ�y��W�U�d����������RS�" PGS���ԝn�n�����O�������~%s��� u�6��F��]��]�����]wX-�^]q����U-�����Z�-Ҡ�b٦���z�q�*��\V��)���V�*x���7ԙQ်�v���{J��_�yIK}���Z�q��}������ u�}�"�>:�q�u�F��*fǶ���>=�76�_iH�O�G�5@�[�md� u�C�7|Qᆚ�����Nyv^��z�bޣ�|��8!� ҡ���H�c㖲�,���iZ����9�m���sꐩO���!<�EŁ�'g}�i��pC�{�D]Xԉ�l�P�~ƶ��hm]՛��?����s���j)����]b�uW�_2G���$  HIDAT�_7�yDӯ��ת������ɪ�j֓�Y�)B5돲��v���+Xf�1����9�k��܀:@]x��^X��)��|�׌�ض��,V����vn�R����N6�t����AV��L�XA���5������!ku��^����|�e��@g��r��$ߑǾ��7>��܀:@]x������{B|�:`66�%6�a�}�}#ޯ��WO���7@���	��u�4�����PG㽧M���P�i\�*
fm��;���ԅ�n�|�gMł�~��@�sͤs|�o>���z���n�:�����:jiw��Q{[v�@mr�+�|��O%�b��P����W|�j8y_Gň� �\����6���`=��xIR��E��|�s�N|��`�H���~�I�H�o�5�Ny���X�@��S���-��	L�FGBz>����P����u׾�Δ�}��L���g��[�/�w��UoԨ�W�����*ԉ�l�Pw��˵���\Wﳬ���h�:���[ʝy!��󴚷��j�!|�����u�NT��9�5��̯iu3y�u���4�� u�'D2��~�%��l�WT���2�W0{gA%���.�L:����Mx����N���7@�[�mԩC���A�g�;՟��oi�ɮ����;PG�C����N6��5u���j��Y*���߿QדQ��{���4��b�u�
�L��;-��Z��ڦҝB"�����kx3u�'h���Շ�Q$J�7����h]
����	� u�'D:��p�ս��q�f(��o�:�Qɗ�?�e�����+F�F�����9T���:F@�P�uZڡ�7T~{�jP���N6�*�y�a�#-ip����������vF!ҡ��������iʚ~��}J^cK�7���5j�ai�%���ʛ�mV���a8�ӯ�~���6@����
uZ���;O���U���~�\�]��u�]¯d���wP�3��2�]fǎ�c�7/co,ϖ�S؂���lz
{e���|eۼ~�yw�t�c@��*-->�KV���6@�x߂`�h�:#Z$@��.`�M#<R:�W�S5P3�]f�6���T.�:Of����>���.��L]����K���lۦ�썥�l���pV:[8;�-]���Z1��|�u���wU��&��_q��s�.��R�6@���	�f�@]����h#	m(Y��F-KBki��=�L\�_���GG��1f=;��àN�u�><�־>-h���e�
؉�kB�@��Pw��%V���-[�􃥴l��-a��pCmn���zj�QaN�w�K��O}��;�T�/�Ҝ�l��u6/i)�<p�Z���:�����:qPgT	u�=ɖr��@�dϱ#U!��� �;s�}��q�SعOE�Q���_m���}������l	�{�6d��N60�D
�=g+5�͘>�͚5�Vs��cW����Jh����	�:��t���F73'%�1�/�Q�C��q#�v�#�}Pg ԝ<q��R�2��4���#�^U�g��5Ch��v�����[�I6��D
����ֲeK֦M8�}���!��#A��T�v��R�m��L������|��d�GY۶m}���=�Ғ��y%�g�n� ��ugOg��d6J��_b�E���ɉ^���\v�s��::1�iN���&=3��xq����ϦGtD��q���6�Y꿥m�u2u�'X�d��^���ظh&�3�����~��ϰ���/}��s���=gs�$���5�j�����.��+�4W���{�N�m�_*�w�'S�>п۸���P���*����0�n���R���g����e׿��/\@���	�V�:+P'�h�j����?�(�y4x`�K�^��� u:B�p��p�NKf������}���ӱ�N�4ԕ%/��f̓��]�u)�}>o��W^��i#L����Z6 �!S���]U�7^?֩c�PGS���K�>c���{��u�W�������+������gP9+C�V�\����<v����i9Z�2u�'�� u�:=��_=����e;���.�/���u����~�}{�E���:���Q};+C]Q�_v޻�: ���;��k�<X@2u�� �� u�:=�h嫣���Y���./�9�Pw��G����	�&��o����'�^'lY���.��I���Q:�ڏ�~�����V��:�����:@�~T��L�0Fk烍��۷S�?u?���rO�:������Fj��)c�ױ��'"��
u�~�����a�cM�xH��e�H��~͆�V�Z��u��J�}4�F����~��Py�gCdCJ���g��Fی!�N��Wi����h����׷�O4�)u��N<$@ֲA$A]�֭���K�	��ʍ-��������}T�$��H�'K �t��M�>�[ߠ�Nq��;��2�)u��N<$@ֲ�P��/U�X�7f���Ά>�${�Ӄ�1�c���j���w�ޘ��~�u���Ĵ�>�E�@�^��D$���^�c۵k��	�����3R�"�Fn�:�P����P��/]�t��^1) �yT:-)`�a����s��s�#����n�
��X=;�âs��?݅u��kJ��`�覞.��U΄�e�:�A�. � uz���/�K��F��,[=�*�{ys�[�������������T�ȅ���ϨG{5��fNLP�>7vm���㋆n�:�P����P��O]��1۹�uufM�Q!�P2tU���S�X�bL��P����ٓl邼��}�+��G��:������Ul��m~UQ����ʧn	x��P�D|��`�� ��zP���R��ӤU���[�>8��^;�-��T����#w����:��D0��M0ڰv�x��� ��l��f��5)��|MPg� u�%X� uփ����XEE�&<x0�>������ݭl���jnՒ�l�+�����������΄8��O�:��Σ�5�8���ꮗ���6�;z���%�]���v����Z6 ��"U��~5�<:s�}V��B=��eزEl��"�6����ݻѰ�f���.��L�N��E� u��HU%�.<PgV��~����_��X���:)^f#�\��Jq+���V�~u�P�w�ٯ�6�F��a2d���ݻ�^�z5��T��:@�Pg��W+)\��p7@�x߂`�h��^�z�o�(�MrN�!S���md� u�:�%�Cd- �0���Ě:dꐩf�:�!=6 ��"U��:@��P���dv���u�[8l��pln��}� ����ǜ��k갦��Ú:#��A�:�@��>`&��1P�]��ՍL�ֆ��:+�)�ԉ��Z6 �a�5RU��W@2u��P'~0����:@]��P�ԉ3@���� � u��J@�P'� u�C(zl ��E�*u�:@�x0ԉ���P���� u��P'~0����:@]��P�ԉ3@���� � u��J@�P'� u�C(zl ��E�*u�:@�x0ԉ���P���� u��P'~0����:@]��P�ԉ3@���� � u��J@�P'� u�C(zl ��E�*u�:@�x0ԉ���P���� u��P'~0����:@]��P�ԉ3@���� � u��J@]tC݁�5l���޺P8�@
�0�p?�`+� ��zP��4����I�l�s�0	P�P�n�&�/+�L��� �.	uO5{��i�FU�v�X�^�T��c4W�fCY�֭k�ϣ�Fԅ�c�
�9w���	� @���.	u��䂺I��:@���nw_��]PWU��Z>z�$MT
��8Xb�U<$@ֲ�.�2u���k��I���>}�b�F򒥛��l ���m ���ye'b��c��ԉvB���ԉ��Z60�ߟ�l�%�CسOf��\*��X�����X˖-[Swp����I�P'�	!@��E����p
P'��L.@�N�B|6@�N<$@ֲ���h�32u�ԉvBP':�C�m@�.Z��ԉvBP':�C�m@�.Z��ԉvBP':�C�m@�.Z��ԉvBP':�C�m�s��.��Y}��F	���fr� u�6J���r68#���_�8�U+�7�4���\,;;�����*//O��&5;�#��d@�/��@�p@��g�3���H����V%�g���y,�K1��1�Vy]&�쇋C���H�}���l ���%��@��u�.fh���b�3��c6�`@����@�p@�,u��M���1� u�m8�/�^@�p@�,uI��MD��l`��0`  �	��P7 f�o1�b,�D�P��:�N�� P' �C5�;{#�$@�N�B�:}(�m ��X�F��D;!�3AЇ"��:��Qk$@�N�B�:}(�m ��X�F��D;!�3AЇ"��:��Qk$@�N�B�:}(�m ��X�F��D;!�3AЇ"��:��Qk$@]�f���/�A�A]@I� Y��:��QO�X�t�K�Z�IM3o�� � P' �� P��4:�i�|@4;�����s�x� 2u��� u�#QG�8e�hn2u��*�E?$6 �	���6 �a��X*�ˊhn2u��;�~Hl ���m ��8%���^47���������L�
�z6 �!�D|���
c
#��LߤXe��� �	�z6 �a��8*�*��y�m@���Kq�	�� u�� �� u?#;��*_&�E��h^�L�b��mq�O��6@�N8 @ֳ��#�cG��&��,�lq�t��zlX�;}�4�������[|�s�%�A��@�R9 f�o�ёE��&��b�Sv	�P�� �y.[��VQQ��� }`������˓��s��2�t���\��u�82�xڤ�I��Q��x!E���܅l���t�N�����P^^��g,�r��V��R���ĸ�{�RQ�a�/���b�c�(]6��^����u : �F�����bÆjVC��ψ~�!����R���$�N�<1mȟ��&����R�״�����k7"���ڠ�~��1��?`���mQXE���9("�-NI��*_��!C>�Ji��r�u�6t@|�����[����ׯ�qk�lq�A��6؂�����+O�枨���b�ٶ8�{��xA����n��iW
F������n���06�������z�֭[�v�4l��U����Ǹ�q۬> �)W�Xy��t�������fp��9��f�N�*�)߉v(2�]W-yS�7_[��{�F��}'�t���}����4A]uu�������Ux��&�� t[�R�B} Vk��v��A�X�%J�����&��*�b��R�"A���6{Ş_��ػ���/juMM�6�����7���gϞ�Ӱ�cZ�����s|v��Y��}s���N���j����Y]]}�����ƍ�zOÊ�74444�n6l������d�8p�o555kjj�}ohhVm555����=p���&�iX444444�[EE�|�QUU���#G��L��Z;x������o߾Ӱhhhhha�vݴi��̭���̎��O����Ϛ��5�ׯ��3[QQ�߰/�nmժU�///�Q^^�!i��ݵ����������oݺu��]+///�}��bm���ԲT,jX    IEND�B`�PK
     ���Z�ȽF �F /   images/c5aba2f5-4dea-4d75-9bc6-8c6f78bbb1f3.png�PNG

   IHDR  u  ,   2T�   	pHYs  \F  \F�CA  ��IDATx�����?��;���۫׽c0��n �%�H`M��������;���H!!B5z5llco������g�?�,\4�H;�>_>be[#i��}z��������y��J(���%����B�*
�
ի�©_rUA_>+#�-9����c���7��S䈢��U�������/>��V�W���ڎ^�O�Z��]�v��v�\m|�&�V8�%�U�חȒ4�4O��������_��(�K�3GĞ8�����L|�o{����m��L�c�J�~�+�Gq��]�Ӽ�ZԚ�<@Y^�j��W-Z��$T�IQ��U޿{�v��$u&��zu��<J�iK�ˑZ`�'Q����?T���9����D��gr���v�N�D�����72������B�Z��L�hiO��ϯ�vU������^�"�$Kx��[��,�C]���Z��H�)���IZ�;Z�P�'�~,��Һ 2�d��Ч52�]�*
t�y��h��He�&&��l���t��^y���j_�BR����P�r;�xY(�36ȏ����N0��P=q��U�)
NWU�EPo�d��SREi]��<�"]Pp*�:Ƙ�	!�/���We���+߅*W /�v���5��ݢ8��e�o�eSą�����y�c�����2�k��/A]���o�]���� ����o���u�qe�3I�P/�"j��8�1�c���p�W��_Ao~���U�B����u/�%�����_�
��s��E�$|���1�c�(��� TѰ�f�*�/%)|�M?��p>�-���U����e��9�1�3�S�&u��ؿ�P���m�{�X6�]9y�BYQ�U|I��c�1�	����EZ{{��ڕoA���T�ǋ+�7�B�j��:kC�CUnP,�-�c�%�8Lkz��h�Y^����������&�]^���N֍��8�1�c�E��JB��gw��P��G�H��8��/�C]C�ʳ��5�h!/|`,u)`t�ڿ����d�t��@�g�.Y��LK6!�hޝ�����^������]���+K"~U��Yn_6)E6o*��l�_�O5X�_�"Ռڱ��<X��S�W�%������������v��/B����6Ԯ������v���U���
������p~����roy�C}����~TN�3t�;�V#�����Vp�Y�`���䣝+���v�3Pq͝-����u[5�V/]m�h|+���) ��H1y��P@B�7~����^��_{�뎵���5(c��I� �7�pwW@q�x_��CJ�P��f����]Z�_�C��1�XZ�i��
�<Ok�W�ٲ��`�ҡk<>�s%T�-���1�X�@	��oyͪ�TI�j}Ӻ6��J�Pw���������;�c��9�������+�ug�_�}Fʅ:}�\k�:!㿹w�1��8��Z�����!���]k{�>�R��j;Z�Ѿ�G�1�c��]8����vW�ӥL�[^�ꋪY��L0�clB���I�ᆚ����4�~ Ș�,�h���-�?P�Rp�X�c�}D@H��nʫ�|��q���|K&0K��+ꮛ����^��1�cl?p�]U�h�Y���-k_�e�P�}c�PT�U�^e�1�;�j�WԬj��e�o0Y2�5��x�P�"2�c�1�V�[^�j֝�ko��bB��c�P��f�TU�1m�c�1ch�ʆ�U�A�u�}�k� ,�.ą���ɷkWx9c�1��e��\Rp��ի?7Q���D��p�jg�?x?]c�1Ƙ	h�잾������~K7�ܸ���+\A����s�c�1f"-�-p�����p����il\Cݗ���"��
���c�1�b�$��?y��6"M�[��ڴog9B���%`�1�K Ԩ�3�Uݴ�����%�]Sq�g4d�;8�1�c,I��6I~���������V����:Z1�<H��c�1�LUU~��돻����H#Iu�7����c�1��8S"����U�N�E��~��d�:��������1�cl	`�,�[Q��۶�DHZ�[^�r�������I�_X��"�L.BΤ,x��pz���2��#���Ggc7vn�Ķ����1�c��l�産f^��O�-Dfn����NGC�C���ܣ]�Ѿ��o� �'�y	!���iW��4�R,)���n嗠��D	I`��8�s�a�qS���U_W;�t�n�k}=m}`�1�ء9\v�=y&?g�-�w�뀷�*��z�⚏�GB4�ݎ7yo<�F��"��P�r���u�).����U'��@Rv�re8q�ǉ����ܸa��R�r��N�6�;����c�}VNq6N��Xu�"dd��/�Ӯw�����߈�oVM3���76��|�=Ha	uW��T-���8�@���6�x�Q8������0���o��I�N������#��zc�1=�-���c���/��Eg�ŻOnƟ��(��z�{ U�EC�ʭ�ֽ���PG��|"��
�`��Ɨn>��J��s*p���Co���?���c�MhG�� |�Ldf&����e��31k�T<qǳx���B��&�1P�_����_�ߺ)(a���p�B{�C�7��K��7����%=�����'�o���hc�16�Д���s8���Il��w��NƜ���7e޻ J6��_���ĭ�H�����+��^���@�F��g_���a<�����_�?�����U0�cAae���K�լ�FϾ�o�Ϋ���W��C��Do�Z��uH1���+'�Z����D.������{.և]���j�{��3����c����)�XqߥzǆP.X���k�������\Q��;��>�bj��r�u^Y�o�N$Mļ��(����sF�v�R�+;�c��ul�7��E��_���*
�zlc�w'�\U}��T�J��P��q�� 6�p;p�][2��A�n�wOݓ��gc������o�{���4r�������a���/!0I�{����iJ&6-�-�����9	���>o���Vu��gb׶�\ώ1�Xڠ�	W��ոk�&��ќ��/�?��ǻ��8��v�U���)��P�0��B���)�&�Q�_��6MT���_����?t�1�Ku}�lT�*C*��Z���%���;	�W�DK6?h��������3%ԉ��gZ�K���T���:�$+ߋ��rn��^0�c��*M��#�Jj�V���N����T��$2�l�K�r,>w�k�[yT�$}:�&��
#.8}���	c�1��h>���X���_����]t5u�yO℆�U_]߲�>XX\�nE���P$xG"˗�8��O��Tu��;�?�Eߔ�1�K5��kaU>RmWv��3p{ï�/!������=ͷt���
u�H�!D��'"���1�|���c��%;�ң���<U��Ѷqg�w�o�r�������C�e�o�H���1��Z��Ӗ/�Kz���1�K�~�pd�y����]��]��# ��P�r���u��[s��d�'B$n�XBo�t@��ӏ��'�1�R�1������f!�0C=#�ޕ*~�}].��)�}T��$u��"�tq��p�c�1�2jT����f��ċΞ����	�&�h�]������1�.�^�V�5�k#t�O���+^d�)3�	��`�1�X*Xt������:��/_����~4
1�\^��$���&#�P@�[P�_kc�1fuӏ�G:��W	w���`��% �3<������B�:-�z�PW���-�C���d2�:�c�G�#ʦ#��l��l|v�9w(�rE��;o۾�2[G
u��7�/	�.��.U ݤ��*�1�&�ʙ������a�B��(F���u�k�[��#	&�B��{3ץǄS�c�-]۫��Kv�_Y���h[����N�
��'��4��tTT��w�r�:�cV6�&�Fˈ��B G��ڵ���
u+�W����I��� Q��I��A?c�1���f ys�/�qM�5��d�Oƽq�*ԅ"�K�@	���O�����c�YY:�������gw��awb�E�*�o%s��sKW���ɝ� �8�Te�[�({�I6����1�g�ݕ��p��`q�j��k֌���C~��o<W@��$
R��ݡ�|!0f�����R�K�O cV���p0Qm�S;k�Ђ�a:�}`RF�/hU�|n�1��C`4=; �(<| *���u��O2N@��Zj�ӄ�u�1�,o�7��-i�/q�B�L�i��6b���N�5 �G|������-=P���c�ڨ�JG�M݉�{!d�%���b�0�]8s���%���f�ZnT$��kXe�1�^:~�M��a�뫗�^��5����<�\!0	〆)wn�ҷ)I'�ﴃ1����M� Gd��6��ķâ��-p�v�~Uկb����Jcڅ�-/��0;c�15Z%���L>��"�'�sEKN�+����W�j��S0�6��'�����Q����c,l~a{Z��m�	%eTtٗ�����������o��H��U�q��a��1�3���L��7~��|e�1�26�����!�q��L��N�Iddd8�Ԯ<�$�o�S�/`�Q � t�%G!�����c��
Z�����̫D����w�ؔ�TՋ`�P�0��B5��̟��8�K $<�8�m�ɋ$�!rP`�KY`�����y�;e�O���vSų�y��A�{������~h�̫f�μ��5I-����6r��=K�Ғ귵d}�������`�Y�lr�����W��wf郆`����(��C��U��\�|�Ud(���ڕ�'�Q?�T!ΰR�����Lٚu�,��'7�1�K54걟?���� ���?����I\8��.ą6�i�X'�ъ�������UU���ӿ2�c�����1_X��UH5�>���O��c�g$�1�	u�u�Gj	� ���N���I�5��%��A�[m`�1�RmoI��ruʍ��e������PsEͷ���r��d=�>�NU�3��t�7�=����o��2o(Z5��͏�1�Kumw��?z��pR�{Om�;WƓ�ڨ�n|B��8��Mx䶧��?N��Q��;��-#A0�c���;�C��5�}�4X]w[/��O�?�I��������8ԭ�_�
��aV�O�i�j���"G}~!��&����?b��N0�c���+~�k9�f�êh��}�>����T T��`��t�q�*���k(������s�tX�;��Ƈ�[��1�K��h�]�+\���(�-�����������a	���]gӭے�p��*�h�@�_�7s����^�����*"a�]� ^�ǻ`�1���p�~�;�_^���e�
�Z�g_��^��Rd�z��<w4R�_^�G�w�ˏ�}�F�}�k����F0�c�ԏ�����EḴ�ض�_�k}.��A��W�x��C�*�8:�>FC��}�_o�ŷ~�܌qy-����Z��iO~aC�cl��P�Ͽ~N��(\p���m��<ho��}��I���.J�C�������� ������3�������9I{\z�<�ӧ�{_�G0�c�uZk���K�sj�V$��v�O����籫��Ѱ�������D?���j��i1��]��^<f
ν�Ԅ��hN�k}G/�L��c�Mt4�m������̫OD~yn��V�R���\-�;�!�Bw����~,=�	`.����闙�N�I_;3��7�X�oЯol���/��r�1Ƙ�Ѵ���:^y�-q�|}{O3K�P�K���o^�D�#��)g%+ԩs�T�Qwp��M��gc��s1��i�|X5�������W�����يH(�c��h�~�t)�R�����;Y(��h�l�Ɩ����G�ׇx��K]��C�Gu4�+�'�}lPeO��~�;�U���E(�+BnI6\.��Nz���h���>t5wc��.�Թa�1�RЮm]�ۏ��_<YnT�)Gqm&�"�(Sk�]���ò>�J�R��0׾�Co�Ӂ*0#��g��i�zٚ�n�/�1�K.2��_����Z��Ǳmڷ����B3�c��U$'���Rc�1�Xb�\Y�*�mk���.)�VM��t�1�cV�
�F���P�@��T�c�1�(*P�}y;��A%��c�1�G���v!P �c�1�0�	�[vUE���W�c���j�;���˙0�c�%����e�����c�1�&I=u�c�1�K�$�-� �`�1�c	�&!o��Ax�1�c,�\�~ �]\{�1��Dֲ�a;��|CQ܈��jz�x��1��D׺9�%�
5	=uB8�c�1�F@$��N�c����*\�**$��WR�CJH��?��P~�v0�c����[n����2+����v!�A��N	��v�H�����Xp�c�1Ƙ)��
&�!or�@°�TdW������-�g�ݛP#`Q�P�c���dLRPqlY��$0O����(9"��ם���C/���Cc�1�b"9T�BѼ0�d����ʥA�
��_n�v$�A��:�c���WPwf �B%�E�1�"v��D�v�^���P�c�1Ch�u�9ؒYM eG���U��O7��gɔá�1�cQ˝�{��8-P͟���G���2�^8�1�c,*Y2j��[��#�Vփe�#�c�7u�1�;$W����z!a+�ò%!�|�w;݃Cc�1��z������䬤dQ�;%�p�!�*0�c�J��Zt�#��S���k��+�Dǡn��"�3o�R(8�o��Z�:&�ZG�1W���E��G	��$���^��z���*���E�WE�a�x��a9�M@;��!��y�c�1�.	�>�N;l�ю��i�A�O~�И?]FѼ�^l8��cw��@hdb��q�c�1��~Q�*���_�	-O���:��HpPB�k��J�Q� ��As�������:�c��Wќ��E��������<(kYn��.ﰣ����"���S杨8�1�c�3h/׼�����pk�c�׏l���nԟ�7����T�['�o�č6��c�1v@�2���z�h(�����ٰ�eʏ	:.�>¡�1�clo�ƓY��.}�]o9�?-OQ��#�R.�V9���P�c����[ 1�!a�ռ�è��c�ug�>��V��S蛘e�8�1�c�3<�z�z6�W�t��F;"
k����P�c�1��!�,cc�4�lT׎V���G�k�ʝ�c��P�c��O���*�(!��PbzǨ�]^}����-��Y�p�c�1��>�ֈ��0a���h����q�c�1�ؾ�u
�
��p�u�z�q�c�1��>�eI�,d0��1��J��"u�1��G$(@d�v���*�
�#�ϫ��#'�'��W¡�1�c��=[ã�����J���T�MXv�l�����P�c����	-�E���a-ԙ+��#�g~�sOc�1���Fvِ]}/mѕY�`�ÜPEC����C����0�P�c����a��p�IAl��J$�!Ђ9xK�ͧ�iӷ��8�1�c�3��.�pX}�)�QuB�O��Ʊ���DA�q������v�w�H%�c�1���տŎI��)��"���K�㏛Y&c�9~�	E	�m�رfb�=c�1���}&�.�[47O������`Z�Z|X�G!�0-��C��]�Dơ�1�c�����hG^}���2f}u=����o���ո˟�$-й�b�����8�1�c�:^q"or$��m�׎.�Q�;B#B��G;Ex�����s�j���w���c�1v@�^	]o;Q|���"���ȩ5��w(� ��%'�:�c�®Wȩ���o�z!�O��`7�������1�cE+K�ucƿ��JM����	6�_	�c���GB��/��4��l��6�?���:�c�Ee�Ɇ֧\�>98��n�C�����F��ل��PG]���dU(z��wd���T�MAߔHH 4$!�/�e�C�v�S�H=^��WFV�w���:�󕜪��Wk�;(�0�i��	�[J�/c�1k�9 o��̊<����px IkioU��K	A��P��e�p�M�.pG*QBmX�i}uk�6�����~j"��f�G��تZw��{�l
�U���7�v���_������/6a���,Y�̈�K�6Oo
چ���-��߆�e�}[����a�\?�J�3���ʐNgt�v����Td+ȟ6���{�mu�w�]����"�1�_�+r���$	DvI�/n�M�f,�� �FF���jӃ/ɮj��*CkK���$4��G�Z���TH��v�G<�=3gfr~�(d�~ˉ/:�� ��_���s��� �'e�v��ul_ٙcO�ػy,o��,0�#�C���������Ù��dQ��l���5���:��)�����-��%���O"�\���26Z�-�~����G�-뀷�z��[z$ZG��DBa�`��f.����G�YZ�{x%�C��fG���Ri���ް�փ��țf~����F$�=��`�'�E?��Z�X�+'���ˎ�L�.}[����{.S����S���� 2K�M�zp�RxN]�ڋ��y����xs穨<!��*s��󭓵O>�|�_p"���el���`p�W���x��W�$Yk���k�5=�S#��T�w�������M����1���Bz0������ZȒ�n��*�N�C�����Bj��:��e�>�ku��:
!E��(?6��ڌ<����4?��P�8��hN'$�|�j"h��m��e�1f=�N/
�lI(�]�@c�ժ��l#�>�p��gGv���Z�U�k!ExD҇~w��ط�v���D.Ԡ�r�v4�������h�u4>]wF@�IK�?Ϗ�/:��Vr�H����ӂț�����S�|_r���ێ�CQ"<���?ZP��o�h��а�}hڥ��7��F�c�Bӧ�j�R��B��R�J��"��fZ�`���AZ�0Y;_�Kƞ�� Z�t�o������.�� �,�k�)EW�#c�&��ޔ���O 㰆Z�DR~L��ϻ�*��t$���~dR�5c������#cR�?��U�IA����E��:R�K�[c�0Hɮ=oU��҇�|A��ն�+qd*�r~ ����Μ�������C+�9��7d�9���F�ΊL[�$6�ћx�����B���}'�s�c�������=hط���^����C�G��64�-��j�n\�(�ηriP�=�9~VS��o&�&��`h|��0��
6�o���vq�F
k��v�k�7c���ڣ�eA}a����G�R¶��)�,��l�qA���`�5�bczVTb$�s�A�`�܉o��C.�$�s�Q�}b��w����cl�(_BV�u�#���:% _OFB���Lo�5,�� 5���w�~���7á.�HF�QAXW�=#�����m�Ao*��7��o���1��Mw�����t���jb�ZvMD�T�ZOPsj>���vc����	^6�GŊ;^3gX�>�T&�lI<\9*J���Mn0�KcblD
-YJ��Esæ�7���ʥ!��"�~�?3��M��5�lh;�x�Ai���v�W��	E�J���iE���d)��z%�B��hGd4�wBn}$��6�5�硺n��������A%�r��]��hBӶ�ѱc;b����w�Y{�
ϯc��tU8+�¾v�u�PU;�����(�#�0�:ѹ����ݝ-1?F钐�Ֆ����ݕ���
�ou��La�x;@ybHr��S��-V�L��x���˜���>�QZ�-Cb�啞������Y���zώ���s�m��e�
z��{��k*��Ʋ3�Z� ��/�����W`ڬ#��ȳ����̿R��/,�/3�����x��?�?T�I�4S0'��w���1�ґ�T�4 �H�5o),>nO�g��nwh!�R�̞��Q{D�Q4,Y4/|�2'Q?g�X��X��o�[t�iߤjyC�z���5#��h+�P��Ү7�/d׆���pM�2ʑ����T�$�PGU�c��{�.e������Oh^s�d��]ki��V�W�z˃�U凇Wk�J�~��T�ŷ�GfED�?h����	�]���0�}�������W��^��i|��۩0�K/�� �Y��_
q'��u���G}LI�d�{�ux�ſa�;�~���at��kn�_K��(څ��agh�þ���u��9�X�����O��{��T�4��Ir��ܺ�CmWe�mzF��q����OD{�m�o��$k��o��⡪�C�b?Mڤչ�[b�.�[�;��(�Te�XJ��~22������wF̬
`����d��t�]0|�Ǔ�e����M2|�$ٰ��������бT��:�hW�X�4>�IŎ�����YZ���q��h�zC	��ŋÆf�;�U}ǌ�֨DU�!M�`�-�4?�RG��׷��:��m}ӺG�c��\9����uC�M�=�ѐfN��+��X�ަ�>��x�:.��g�P�V��ͭ�Y2iō��P�
���!��V���[��|��D�3jg������ds)�z�Pv�ٗ���6�Z{�n~��q���1�:�y���}����ww(<�ew�� �@�7-�w�m�Ù��e��Y޴Hj�:��F�AFt���`�}��B���rg��G�������ȷ]��?J��N������l�ȧ�<�А��,^�m-��ɫ����0�5�u�`m.	!���)A�ժ�zK�?M��Iy-�F�N�Xl<Ŵ��/�9NDq�9�Zz!v�o���@��dW����X�}dWF�x��࠺�W�o]�*�pG㺻�~�*�/���?y�lL@�
uFW��J����n�	�����5�s�=�z��
F:���d<_Z���ȳ`�f�Y<��=QC��]�7o�c��3�X/�����ŧ��������c���,�\������ ��{̾_���%L�}��M�y�G�^m��Q�F��j�E�<��^��v�F���X�	h�����[+�	�l70y�S(�ꌮ����of�y3*5���+g}��Q�̍X:�uvv"+++�3:�G6����?)��@� 
�KU�{݈�i��t�;g�����KE8}���K�3�7z?�C	��-�0��[�Vd��uّ�˅�Uzޱ�mk��B�+�X��`�]�P��"A��[�7̌~h-ֽ��ơ:tf�e�U���e��Q�̶P����z����D+)*v��
��՟��bR	��X�rfkk�Q����ihi|/�cbii��h�;�����a����e���vln-'6�H�s܉j�[��oZ���vs�w���+ �=&�%��q�Ǝ��@�k$��<��g�1'-�Hnc!'�푑P�Ȉ!�9T}�T�hμo�x�����D�-M/�tV�Y��:�9,�c�!C%gC/�v�࠭	�K�r �P'�X��0�2��YYQ��Nr�x�K�@��"	*�Es�!�h{C�ksk{#>	J�0�x@�_����i�Bu�!q#s�(W��~"�����d3�"�nM����j�[�+��/c�1��NF�l���������1���>����}���H�SiD��k���&ja�	 �Qd����@=�jD���Q�p8�#�m��'2VpR��S�1�Qh�%�g�˅��L��Tf�DU8Lm��� ��Q�1v���	)J*�04g����S	j74���+O��ػʴ��%d�9&�V�J��2����@7
�*`���݆n��6a�黳Hv���R��N�H$�ёAӫ1�A��Q,�b��G�.J�{�E����y]ي��r�y�lQ��АMu�O��,S
/�]��浯�$�u�%�e�������BNpH��>��ȉu;�>2�㯌1�.TU <j�#3���ڣ�S��\:�G�!��/uLD|FJ�yKչW�n��E���0��c;+��X�ap��oT�.�/�a`���)at�k��vմPgό\�Uilug�?�9��-�~�AӶ�1k�R����w�n6v̐�C]YY9$铟���AD��a��Ʉ����w�3Vx+�/�'�����a���d�����O�;�.t���U��1�D�!��PG�١�v���h6tL ��WBfF��75,�����?�I2J��2��>k��E�|�%�O��NiGo�|u���f�6���ڢ��K�ND����[B����'��VS��o~�ED�_�7I��o�ۛ��rs�xǾ�z�#�\��?"�L��C�#3��!�96�G�+ZX=�J<Fv�R��3v�Tq�4[h8��������`�޲�o����>%(;�����γP�鋵�Վ�,�>P�O�`�K��4ԭ�[�q/�X^{��E3C��䠗��m�)Q���v�Y��V�V.9�<�M��y�cnͥ(�S�(�s�#<*��En7�	����e��F��/���y㟆���B�u������/{�W�ؿ%f%�w�3>��:`Y��A����i���F!F��=��W^x�-[n���\�M�>o������a҂�7�ř�ǆ�uߢ��*������߽�s�}�@	�PO��G��W3R̗�v��s����wg��������՟8��J��V;bݼ Ы$��4P�����z�Ѹ��U�<qBAc�M�g�6�g�16.�}���z�m�� �\�ӂh��ӏ�
�}�"�ͱw0P�S"�P���i�E�lPW���u�1>��z��=58�����C}N	�3�����vC陔Dć��+�������~�{!.�M�[[}J�z#]�{�m�}~�����,66��ֆ'��di?H�����"�'�Ǯ>v�%�1���5is#{����<���e�<���S�ރ�����m�=��A�o��7�XoY�ID��ۗK+K�l^�_F�]Q�¥82�;3��X�7��b�Q��_��M����>{b�\��BL�{n\qG�-u�e�ߙ���Q{Z��X���_r��lGɢ��r?*^~�v��υ��s�!�g����~��Q	����1��M�C�Ҩ�@,>��t��^��{���F�Ȟ�+��e=��C���~Y@�xɹ�7̵����h[�t�㮨��X{^�Κ�3<����H��7[Eԩ��QC-6��;i
v�C�q��w��xw���ϐş�6�?o۾��"�V�E=���^0;��dqH�Z����"}�ȭ7>՜&���l҇bk��V�~��x��'��M�����W�KS�n'F;��k�TU�[�=��������v�A�}�#z�����^��G��N�k��_�FW�R'L�1!�O�|n�+�eW8V�V���w��x%Υ�79"ꙮ�Es'/�s�b����:Tugu��Bv����.��g��h�������n��~D��]yaoV���*9��6BC�ޫh��N�N��T�{p�[�����3*kfaRI������	k��v���Q/[B�ܱ
�H����:���MHf,��T�?�Ƃ���sb[��۳�|x=�Yy������*}/Wz�F�!�=����l�E6�[��G����2z�t����c{.�
�����B�hy�_W��~Hk�G���y��
T&M�ѩH=�C��*%f�������b/���(����Y�3ar5���cU�M@K���w�hn���Ƈ��_a�~�Zc¡��qURbhÛ	ihh���`ƍ��1�=�ѣ=F���y�K ]��YT�S���Ε ���~��lu��;���9T:_7���p���K{�eC;.$�`�؛�L�^v!�N�#Ӥw����7|߇vd��6e�1fQ�Zh�&��z�/-.�����?�D֗eC+��:|F;�Q�no�P$ ���S����mi6*A��O�Ƕ#h��´���Gr̨�L���g�1�8��5?AðXi�?8(��������~[�r�� ����?o��7�n-�#C=X��aTB��n=p&��N���\j��E�t����f�1�p��vt��D����A^���ƿ����Q9��%�%������W��v=1�Uv��ë��M��M��1ڕ�Ɋ��v�ŗ�֮3�
��t��Z�3c�%ǮW�z���v3P�ٮ_b��S��|і`�:���ͣ� ZU\�vh/4U~��C/p���J2�|ɩ���#��|��Q;��&t�16Q������P�`\��A�b��d%�v�͏Q�X3��|��ꉻ_����EA��x+_���s�H�ʕ��O�OHt���c�k*]���k����G�4
E(���Q�W~�ۻ��0�n�as�3��|څа��J�oꩢ!H�[�4���>9v���'�|�TK��n���)KEw���˝Ԟ�+'�T�lhy��?>s��U/ZZ�=# w^�ϗ�Li��a?ϡ�5І�����W�:��O�}��B]�D�h�ǵ��;*���@ޫ���cG^�6�k�0�Ψ���.���LB�����/W����ڤ���=-��*=8��dkL�;$��P�٦�xQ�(��E�
�ε?�4�lI,|�m��~���X��D���Q:*[�ƨ���2��e��^��\���_߷ k~/UU�3��w4���F!g�}}jP�a�T�
�k��
���ٰ��(;2�I��	鵣]�ڞqb�}���S�-��������pN6:
h�Z����]��g�1������h�Ks̨�C�K;_�_���a�Q$�*cG�X�z�c�AUv��B�{Z{�(���S:W���з�nZaa3�A-d>���w�V���2��Z���w�=%��LH�9g�����S#ȟFf�b(�P6����^BE�p�D�Ev����y�2��ͪ0v��Lz�Վ^:�vk���2��C�z%�����5jdd������u��\�]/9��(�_�����G��>ni!���P"͵���|;�2�P���Z�H�K��U��$�_�Ơ{7��M���(p�)pd��9U���/9$�7#uy�����j/,}R��>�Ѕ�Pt��
\�*�Y�>�K���B;O|�c筦�)Y$W0�:ul�Y��BϤ�m'��-E�16��T��M���Q���W��\6��/R�fRi�fP�K�����>�/�4�cO��t�=o�zް{>9_%2�V�Γ��Qod�H�`1�O��gP�W����("Y�K� N`��4��D@�����c�I���1�cl�8�1�c��u�1�ci�Cc�1�X�P�c�1�8�1�c��u�%�;���O���!_-��0徧Y�U.��9d$��u�BPկ;�.�瀷����'A6�SJD
#��*TU��q�RH�cq�a�������C$���>���L�����r<?�K����~�[�M��GG1vf}%cl?޾�>x3�����Ŝ�#1��s��iC H�>00 ��s�۟��L�z�,}������倂��I���&Ams!�3��R�i��\XX� ��;W�d�Cc,.�]}@�~�73��hl֯���C�:���n������Tsx[��D}����Y��P�c,���!��z{9�3�	u�1��~؄���w~؉L��S0��	upxT}�]��>m���H�Mu�������^�+%D`,�IB�����~$�߃�����[�B#��@�Iy,�H@u�F?N6j����=��Q�������Jv�h��(��<ߤ�:w���J�2<
����B�ȁ~_���v���7[�q�)���|3�|�������0�e�m���/��c����
�0�;j�D:�67�Jk����_W���O������R{4ܮ]�6);Z2����\��P;�lE�X�4:7���c窟oۄ�:ɩ�pV3�Ș�o:&��.

�F@��[l����@��Ч�d�9��Y��-��|�zm�R4'���o�o��ϗ1Ƙ5��@��0�g��ɏ�=��T�KTxKL��*�v����%�����Ύh��;/�'jsk�ZJ�|��D��3���ѡw(�*�C��EA͏�o�xЧ��:Y��$t��D��vK����]��7�� �E���S+��ѱA;�-��c���EZ{��2j��A�	��#����Q���Z�������%ǃ�g�F��Vv���`���7�>�\�_u|�L�/�n�͵��i��[��*�e~�O��i�xNm���{��|S�MJ��t�;��aT�=����S���� �ZmZ{�Fpp|�R�u+?&g�~x�eԟ'c�Ɏ�g\�N;bJ���[~tH��L4�0�~�|ɉ�o��Q$FI=�2:_v����E56�zA%v=��KG�#Wur ��_�/�Zk��<���ѷe|z�l.�'�7%��S��
-O��Q�T���{UL9/�ONL
U�K�z�]����$��B�����zޜ��Η>-�>��v�1���V��ם����Bd��Z�?Ɂ�/��:=ȕ������=�����(�'߉]�:auq�:za��H��7Z\@$�uCI�S�a�)���խ�p���6>솚��c�b(�M���DLw�F�a�-O&�c�:��|.����C����#ǆ���$w���(\ԟG�y|ώ��՜@����`фL��0^�n��������wR{(��ByN�~}dd�16�83��#G����4�O� m�r%�q(gԏS��[�ܱ*4�Ϊb
u4H�.ڥÉ�7-��>�.��\�����>Z�ADw<o�7V����(��h?Wc�y|/���m�:�\c�`h�'�D,Ћ����:_OL�K+zi�̑a��֫q�~ךs�c
u���:�,ŋB���*f+;&o���;i���.����M�����'�|�sk}�c,>U'�.�V�[�$4Vķ���n5'�m�ׁThh���n�U�0���d=�Z�yӊ��镱͒U!k*���9)��w�n�D�cѣ�3���(�)[sJ�~�ѷ�4�#�)VVC���Xd��I��o��PG�N�N4g�R�����W�^%�Q2�-;:��u3�ҧ"a�{�f�##3����#�P�G��Uh�۽��c�V�V.5���nw"Û�~��;)�V�6m�o�Ǚs��%g�'����]T�C��]��X��6�+C��pND_R+*�׳с�f�n_�x��"T�Os�u�e���rA��ثC��(]oioԁ��X�v_�̣�j!n���P]7��eڛ蓮�H$�ݝ-h���mـH8�7o�0?���9��c,~��q�t��)���G��f6�
J�w/
�?������E�c�+>,��5�����,�cE�2����P����=���rk�vޓ���ꭈ��?E�ʛ��^�Ѡۭe�B{�G�תxalî���e'z�s<�(��l��e��c��WK�-�cvm�����������S�8��'�,3-b?_����ȳ0{�RH6�n�@Y���H�톗����^��y������f�16�]E��b�typ���bڬ%�t,���p��z�~Y��l���_����6�ڟ�o��v��u����j����v������DV��7?<u׫����s�аQ��T�=O+կ�:��N��ç�Nd���#��Wַ��׃�v�(h����c��p�`���S�nap�Xތ�_T�Jϴ�4�əY��8m��'�Ҩ�q{2q�I_BE�<��o�^<#r��{W��ޤM�c�ɮ��Ӕ���/�i�\��KQC#L'�q)�+��g���1ڇu��.}�3V4��޵��64����}���[�;�m�<��Rܣ�屆��W�̗n�8.d3:�h~����[u��erfpP�;��8���[69�Ζ��Jq㖦�x���@���Q�U,��k�q�L�盙��e����X�MY ������E6�nS{f��1���c�%KuF�j�����w�b���^���T�v���:Ez��F���E+Q?|Ƚ5ĩZ�k3p���i�/����x�����|;"ή�`���(�z�	!��Xȡ�����a霻��
t{�������e啊cB��7�g1�PG��k��/��r��1�=ʫ���c����=`�̪ �:�3�jp�`�����!�U`,�8�.�zvĆn��)����omx��q4O-�PG��=K�D��~�����	t[߲��+p��܅�Ǌ[�K��S*�e�ˆ'v����ͻZ־�8�x��U�Ϋ����$�o��L�?1Ĳ�:�����=�$N��f�;V������1�P���X<�4|N���^�vF��^1�J�tJ1�����x)0��˝��A��6r� ����y�9�E�<���OC�������1�ZfЇ1cx)�+�W�=h�#�W�@�q���O\��?ʭ��72�*K{�Իg��â
u�����r@��m���j�/т�W�n��z�)�U�CC�c)��Yn����tc�a��K������C�.���&Xr�~sK��ݕ�ڊ�L��P�Ό}�ۍ��l��"y&�������9ǚ���d�aG��=�˨���Td)1���4ͫw����M��	"��7�W�̉��W�+WA���G�<�z�n�C�[?��7��+�V��۝��7 ԅK�����uSӂ����J+�蟴��>ƙ#k��1�҄3�X3:u�z]T3�L������M�o,���n=�;hQ�`�_n�u�*i��WY�A�;eB���&��͒���0QX�l���hn���ؖ���}R����D�����w�����l�U�fl����;8YN����N7�YD�g �{�yjԤ���#���U՘�Qo]E�tl��F�����j��+�X��`��z�)>�����uѿ_c�f�*��3�=Y�����D���{�o麩�Z��I�C�c�0��V8��PXdl���e�7�XfW·�76D��cRn�ok���k66�TUX���R(B�op�9e�����f���}b���Ʉ�9����V�8e7�[ˣ���Ɂ�B��i��/���Q��GFB],�/���UѢ2"�>��ט���������k�Z��������:D�mf���GE+ �4S3�Pg����4�����"�Y�����Pǒ�Ց|4�O��"�|۱�dc�s��%5�G�_��΃�>�؊���Q����bS����L��ã�9��fpg%*�E[Q&Bf����C��;���Ru ��0҉d��Ç�k���=�UO�Ƌ�DC��W�0[?WCH$)1+N����`�W��;?��#�?6�E
{�>�(�@QW5Kg�Q�~�V�~�5��UH�k�;ҁĲ���6[MH��~;�i�{�.ѾW�v�	���J	�c营�Q�hnԟ�T�~�R��t�D,�b���ѷ�k߿L@o}�1�c,P�W#¡��!ό��0���?�`I.��>֊�o2@�#�m8@ۡ��X����Ъ���KW��Z�J68\9��P�T�|t{�u���f��3�:�!�Q�c�B��zK��@���`�M�Q�����,%4ֱm&���^���!W��*p�U�$nj�!Q��Ѐ��@��,�dw��B9��$Ro�Y�AC��C��â�j
qw�ܞ�Pױ�CC��$���]�^/+�z�{Q�(��Z���+�����AHx�����%"��2����Q�dxT��}��*W��o�����-0��R�ͪ0�'��HYT�.�o��4�Y	��et��\C�� Wd�[苭�j�)�ظ��_t
���i?D��}�[�X�%�������k����$0B�K&���A������[_ǴYKL}}���6�!�[�	jyÙ���O��o��+�՛`����ծ\c�c��)�F;%̌�N3&�Ȫ��z���ii0�tY�w���kt"�hWl/2�o���o�׻m-�L���[OCQ��^u�1�N����"��=���jEQ�y��}�)chy������Y�y��F�.����v��h��qj�]��h^�0#�ЂO
���ƿ9UKC�]�;/�^}�}�kbm����(��h���4���En����p���?���)���_�L{�mz�9CǄ}6��y��1�҉��f:�g�9^�o����fl۲��1�n[�s�h������|����E��.W��M1n4�f� I bҸ_�ͽ�r�$@ʗ�
8��0c��{S�K[f�7g�l˲�ygg��|��M��wf睝���yO��A�����s�G��>�5';S,]L�oMR���k�)j���u�.�"�D*=Sˌ�K���4<!_�/j�П�gM�ۓӯ�%����&��J�c�@{���Vl��4.��V�D�$y�{�*���{�2�L5�S�a���G������p�a���Շ��eX�$5�Tjw0�5��dE�:wq��,��j�T�Z^��һl���˅�%��L��*z*������,ȺP�FH�Y~���/4�t�������^��~u��f��%׸��'��~�8�Rd�!3r��͗�f�6]�M)�׍7^~]�\{���=�0�D���v q�XI�}��Uz�/Xx��������=��>� ��#ڝ*!?�UfF��b1ȤO����C�&u9��\{P}���ӿ�j�1�Rz�g�9FLoPvr8���g�~Ќ����*c�[b`e͆Ю��߽�����pg����M��O���>p�~]-ṝI�e-� 꽦e���6\��p�īޏ���}����&u��툞��a�я�
'f@�W���W��Ղ%���]}-զ�2����0��Q�La7�o�/.�܋���o7n��_/����U>�a���\T��<��
V��-Nq��[c��?:���J���:��2K��5ō�v�첼���{�K���`��먧�7���3��!\��-����~ͫ��[�O�7��EӍUWsk��c�=��:{�⎒,()��|�.�!��8�}�c=�a���ǌ�j���Q��h�;���+Y�v��˯�s��"���@ku����Ǖ4��غ�<�dA"u�	��-;,�|�z�V���!z�,�Sm]M���9T�`hel^���ܹ	��K��1_=r�4}lC�,���^R���E�/���o2���b���7���s�+`K�*eD�I�5t!/]W�>^��m%]�h��%ɍ���][�@zf�2
��$RP�ޞ647T(OQ���4���
sd��1:a6��թ�.M��j��/�a��e��>M�<�~l}��
22���ؘ8���J�Z!��vT�8�KG�+=h�Њ�nhi�a�	!�"�B�.�o4]@�0|F�>d9B�Έ�	����6c�)z��!���6@V��:?�z[*N�h�95���n�U��K�#��[H��qNA%{��HP����t� �ǚSz���n7�}�,�9��K=^)��@/&g�r�aN��݄�}���n��$�7��b�j7��]��:5�A�d�ۧ��7�>�~S�yS�]Z�[�H*	e����OO
z�"�:Jov�F�|�[�S}�3A�5��.�ߣ���٥:��a�IL�V$�a��@��0i�i��M�ز��6���[�������s�[��R��3?��i��_�f�U3�-�xŁY_�)�j�Ҳk�&^jc�9S�{e��ގ�7�a���|4�������6��5;���ִ�)șҼ#��	hr���~ӆ╞pJ���o@�K%:вs��v��Dō�s�Bs�#j�2�0��@�	���Q�£)�Lo(L��-fQ���lȻ8:�SۊW��o�h^��:2����R��X�,�^�C��ItW���`C��	��wp�T �a�9��8`��aC�҉:�`({��@d�Q�.��`x��:@$�o���7������;Vp�wB<vTv�L8��s�b�B~
���}pH�Q�/�0s�BI|�<���#�C+Y�A��6�$#�O�c�<t4_�/zv�v�A�#����l�;�cS��MV�㫮�V�4`G��^��a��KŔ+�;"�d�a&��"�Qx�W��V�Вhիv�S7�4m��+����q��6`Uoڣ�C7�.ݨ.͡8Qx�qy
lB~)@��2'jM��Ό�O�Px����J�ͱm��[��F���a�IFw��ڌ(�ʃج�E*�Ѳժܝ(�K-�\�|��������h�؂��V��'/tTt�-Ek�G��#y�9˼����\	���;mZ�J�ؤi~�5�5.�m2*u�\����0ÜZ
=��ɳe���KV�zkM���/-CN4t���D��KY%�4�~��_׽a(�h��r��;D�g��҇�Y�4�h�Fz*�H��Cƹ������@��|�C�0�0cA��(���I?�[B��(8�G���G���~�Ӟ6Ǐ�>Xc���Iݤ(�x2�.�Lؾ׬l1Y$O�+�)�.8�x]M&�Tޠ��H��~��l1�A$��!.�@���Ρ��V��A��9�aF��H�vm�e{�PV�(,ʞ�ΛEK�TwN��G���G�=��^T��E�s\n I��������d�]���8A����;�6����#�%&�0�g���i��.#��I[�m��(o�E�%�H;>_�Šw��,�ȍ��0)�3�0�(�>�O�,ٔ���oH�Ed�Aa����z���'��Zѳ����`K*?S� j���5(Y���-�ߩ�qQw"~Y��LQ��	�ð��a�a&���Θ�*y���93�;ĸ�:�a�a&2��c�a����c�a����c�a����c�a����c�a����c�a����c�a����c�a����c�a����c�a�����3[5إ��R��SCa���6y:����f�	�|�9��0�0��(�+٣��'��-2��������N%��l�|�1dC��86�ny���5_"��h!�0��<y���T.�� q�j5��΄�3�&�衛(��|�ɣϗ��̈́��O��lD(�a�	2	E����T�/F�1AY���WoFO�I�œ	�,T��ol���Ш�����W�=�f�O������:3�HH��٦^��M�P��%YM�~������V�Ò>߇��~����K7alv@ٲh�=��m���D�|�a��đ6h������54萐��E���(�#3��Y�K��̠��z��/4_�&��e�Y"��n��jF�AsT�w4tu����TBR��'��K);�<Zw[м=�n.k|���%M�i��E�by��K�|[��o�0Ì9Sr�z�A{dO���E����e��;-58R�]&!�@�����_*څ��5Zw[
bR����o "�H0D��g�u�|�Sf�Q����J'r�f�+�������}�Rf����Si�0Ü��e.��6ɧ��7&G�K�H9KB�;ve�r"!�AΏ���.Δ�1;C��M9[�o��?���tQF�^�Q\���<c%�yжۂ��lN���7��J�nO�a���Z�����h���$�a��L�9y(����|��
4W�".%箜��x��!��B�Jb�"oh�l�n�����w"�X�D�%�H�Hb�M.4~lE��aĻ�-��]9�z,1�7[r+S��#5�����<Ior�|S[c���M��Sn抗��z'�Z?�0�db��%��ˋ���&�"�2�q��.�t<�E]L�l��(���b��R�Pūv�����J�a�5e�nܐ�K����V�a�G�a�:��JeAg�M�|���c�g]8��c\�
��A�)����3nt����a�L��J�u%�	e�N�������Nq�ū<JE�� i%A��
�%�V4�:
�,��[t�P�u�|c=ǎ@��N���\�4ߣ�90Y�s�a&�^ލ����ϝ]�[*۱����DBٞ)膠���zQ��=��A1YA�t˂
�\���\vѺ��Q�r�N������T��"W/�P�`4�D�^T���7�af
��Эl'���P�Л�1!�^7�nZ1˻ث$�E��/��5�%e�/�L�G�4�:ZO/�ܫ\�h"y���>%�@o
Vx���h"i�i���;�a��,��-��5�!���d�kB�Q}]iTe����q AY������w y�_)��P
rO�R�~˒��N*�[�Eo�	��0��bB����(ICL�&��e/^����z�t�A�b频�˼J����ޙ�x���h��[�{p�Ψk� $�h�5W�Bi�����3 (ߟ&kHI����p�zqyyQ�>���k���>�ш��,��'�d2�'y��݊ޞ���K�zr/��i��0�����;+�s��Gԙ�Ad/�.d��R��$�l���FOW+��:�;����I�yS�eIk|��?_Jj�t ��A�T��R.,�[J]��6E�2���˘�Sj�i���D]}5�����uY��˗������<[\���R���y~�V�'� Z�w�f���U�%3�gͻy�g�b�ƻ\��,ۅ�7jx�������˰���H�");���~_��=#�eLK��|����~ ���_�N�X�'K��U1�X)q�9�u�������z�3��^������Tq�ĥ���Y�?l�A>F֌�ƻ��>�p�IbV���c��z$t7�8���X��^�:<�ku�'��=a�<����c�H/I��z�K���_{��hzi"̖�עK>/w��k���&_��ѯ�T����ކ���q}݌ްJy����9ː�?f�H{��ׅ��;p`�&�wC��|h�n�ET��z�z5����4ھ���3����F�?u)z�"GJ���R���y>�Y�����]H��S�X��#��~� �P���[c~�`����ʟ��f�����~f�����~-{�Ϩ�:v�>T�����L�%����D,����bn4��x�=�b僶_v�?|)�)s�h~��u�Đ=+	�o�y���./��ϏF����ٰ�7&��t5�چ�ɚ�,k��cuz���>6��Kd�rܠ�Y_���Ռx�˾>gؒ؆���aǰ1�fb�U��~o>҅�~�w��݄��^lv��;dQ:\��^���xCTnm��;4��*B��c��P���W3��b�q��:�|i��!�6C�C|�ϣ(��iؘe_�)���t^t~Cd�NƢ/�����|���}��+�_�&���}�5��䝕}L�In	����G��A	����A$��f��p���#+�t�q�qI�w�
�}��ؽ�-�����E�>�,E��
*'���D�j�߶y�L�B�XS�ȩ�N���w����m�����i�W�;�`g)�ލo�jQ�2S�Q���&T�b��׬�zx�X��P�f�?_������̯ʓa,��X�Wn
�ZI��Y�|�3q�5w��U�)׹.CVn)�x�1�]}B��+���?��6�a���������EŎD��b�&�Un�L,_y;�V�"�d���W*��W��$�!š�m�UK���48t�+̨zݺ?�5\�x���c���'U�nY����&㺢��q�Y�)��n�b��c�E��<�lD��}��a��+j� ��<��v�����ٷ̼�SJ�B�(�Ç�mVh%e��SQjzV~�۰X�����|���.������u�ޏ�6���ܧ^H2�0��$��x]*wF^���.Jv�4\q͝J��s��뾁W_�-�~���Vג��ѶWcH�a0!SZn�x����n���
���y��Ֆ�ϗ����:O��
!�@
��<!P��m�+sf�e��=@�z{[��ԟ+tC��ꡖo�~��fCp����(cU��#]\��|�V._u�fA7�^��xk�����cQ�0i7+�5YL�OԡȖ��`M9Θx,�����YEXtэxo�SB�%�!ꨡ�h�4�xQ������g�p�AM�k�Qq��߯h� �q�RIH<$�&����TA�b�6�{�w��~�a�����i�������&D-�Ԡ�\��}X�<_ѵ�s�Bl\2���d���Cu���X0قx�'`�af�Q��A�/�4Y��s����}=G�x��� 43�^���[��X�z�ج���KK;�x%[jߵ��R��kjޅ0x�槻�n�����_9�՟iZ.EA�U�.V�k%��~�����_�<^��sw���ބ"�\��.plf =��O*��b�%<�:{	�d�«�D���=M�@}�Uid��Bt6vc��?�%�-��ߺ���Q��>b�gOu	I�(��@�30(���~�~�Ǎb�E��c"�Z��4?���a]�u������{��dA%f�LJ ����kW�x�Ib"����Q�06��z����8Rԟբ�1G��|Kf����dRRs����:����~ r�-�0g<SG޺���&����"�_���6t��^�h�����g](?�����7]Y��egO�&�l�z��AS��Љ���.���[zH$I�!�wx�guA��Ƚ5&�창	B��՘��S}���� ��-:_�0�����D�%.:+�3�Lrfd����8�o3��*�Xhu�x�x���#�r��>P��=QC�����uƶ�
�G�c(�l_����꯽�n��D�Y0���a*��x:������"���v��-ݒ���H���z�
S�0�D��8�e4CJl�����l	��C�B)ZC��HeD<]��A]��*.����y1�Տ)JJՍ-���#��a%G���@iG�E�Uۧ�,��gd�N)VO��E���ُ�C[1�ǲ�t���F�`��iĸ��:űB���y��?������g=������c�������;�X��O�!˩�+d�Q�b܈1�y�z�2'_W��y�3�x��0N�*�f;隙��?7!0�ELp;���?�嵌�Q=6�C�P�!��Ȥ����*f��t�	:�K�T�^oآ�	�����<=ńB�y�1sK4�e���;BEE/~t�>d&�8\��OZܰ�I���i�i�ׂ'�g�8O�p�A���1')y�ԯwR"�'����q���^v�|쓏e���n���D�cx|]�aǎ�������D��9:N�c���s���Л�7bl�$��M�6�{�u��?��׌��tc���/�u���^=.�u�И"g�b��w��Qd􆨎��;��#Ei�j]��uju �dA&Hn��|��u!x<�p8�7��
v���L�񧽳;��?��W:u{�=��l>��=�{OG��cy�#3��TT���x����S��ν��~��٩��ݱ����ޑ�9�?0��{�g���A��qa��~���y��{k66�De��h�8�CS3N��CGa�_�i�Y�a����Z�{;:����}����ӷH��=q쩮+�!�.�ׅ`0 ���ga��b�s@C���`gNZ�5b��*1� T�,(^y&"����bn`[r`�ws���U�����+ܚqw�=)(&�<ڤ�_��*����G������Qh��0�B��t�D���DOk[����5|�}טcj��m4� >غs�c�W�(�X::v���Gʡ��{�9f���;4��w(�j���L��<��U~>�A�+Z��sW���5*�"B(ht2�t�P���$��s�ڛ B�aȆ�#Im�0��`��Ǡ�L7��7J~�gO��x�����j�n#,1�3+�������N�ee\�K(X�ӭ�"�~V�����#JK�i�;,4���X
�a�3����//V~6����KȈW��iAT�>�{ݚ�>��Q�G�u����-�-$A'�aKPi���^���s�T�\�*в8���.��銎�2U*��i*@�<ˏ�����Q��d������tj��^zs��Ϸ��v��p�F��Ԟ�V�4U�#���c��Jx�LB��衭8�m��t�4U�6I�ۧ�S�S�KLԥ������k򏺈��⳦��]�X1�ߤu�&��QS��4=��k��V����&��*s�g��>G�*��6O�|� c��m�>k!�b׶7 �M��EG�9fr
EG351�c�J�^ލ�O�":c[*��-���Y��~-����U��_t�n�k��Bヲ&s�h��M&$��G����w���?;aRJ�����S$��Vq�O"Q�W'~�9K��5��+�������$�	������<��&N+���0RiM��W/~3n}�
g�0�T_��Cۄ��zM�'�E	3�����V2�4��v$%%a2��Эl'����-��p���W�p�s�ʙ�5��iU�QWsPhW�	����Hl��˼�CO9��5��%�h�� 4rG��Rf{~%����}_	U�N�5*�ը��Z�uY|�'�|��Y�B��r��:�q�X�^�%�p�]�})�7`P�|1���X����g\}�7ê��ׅo��^��z����a��E�1��o�%V�=��i�Ʒ��+��$�JWg36�#��.�6�l�i�D�rϼ�7lY}��ϯٱFXR~�����t�܋�g{*�'�I��P?Wg�X�q|~ %���*_�~�M�?��Ꟍ��	w�ޓz���l�S|9��7:��DA���?�Wf���Uow^{�Q�z���bQ�0�'?=�v�n���g�'2���N$�+)R]���;.^q+�&�U������QH^�"��<��@L����S�������^|��U�R�����{��e�^/��7�$��eBg�$u-�Z$At�	�~̼9xv����w����'=2Z���Y8�Ͽ%���(��a�����v�b�|S�.� ��u����?�ŗߊ���{�P~d������p�X��9�aF?3��3�K�}$��Q�[���J���+���}��ڿ��"�~��q�Z��-��Y�1�'\�7�l���%Uoَ�.���.��Wk>x�I|#������ϓ���D24D0u5k.�	T+�ݦ\��o�#5�����]e���������!�Fk�@{�hJ��B؂����ɘ/9E3]O�i����d�^Z���y�x` ���=�K����ː�]r��`�߇ڪ}ط�]�6Wk>����c��;dqeP6���8�s�˄�#V$���m-5x��GP:�<̚���ly�>���{�w�t�k�CH9Vz�_O��^@�`,=��Y��;X���guѽ�!dxG~�ꍁ@g�Y��O'�HWf,�[e!��<�+ټ-��ꉐ{�e�)g�`��㌞0�g�i��⭮�T����ml�E�I�/w�����&�S�-ۭ��7khGHO;�e;��fw*^�ظ$��6��7==���!��&%u�7Xa�����0��K�a���T>~IE-��H,���b��2q�����p�!5=1���=�*��
�=�q�@�t��Y�PꇖJa�U쐷d߀�k�V��|}�u`��`O�z#� �8l�\:-R�:�ˀ��Ȼ$�~f������t2�F]�1�l�!�;����i(�}^��5��;!�����e��:l{i7B�a��b6R��F��&)�ik��8&�Z��#z.R��ۭ�^����>
�*�Q��~���R�+2��N�%\$�{�Ƃ�\�D����j�k�����<4}`�]5��3#�Ԥ$}D�[�n7�)���a�QGgc7�\�Yٲ��+�n��Y��#�
R������R�6(��9���HвM���>��)�߳B����дՂ����m�IkٴH",�h��u;f�-Y����ڌ�(�+O�Z��/��R�#M_�MG�S�0�T���U�^t#rfd*o��H�NT�=�8W���"eܞ�b�,�:>)Z��U��l�>��=���Yq��y�*��1��p�f$i?`A���LN�tV�~�_r`�gܚ�����aD��6��������7V���a�8�4+۫�߀��Y���f!1spل�z�]��K�p�{�x]M=a���ǈ�W��iw�1�z0�lD�[��&{W%��k=��X#�c�ݠ�2��h���F�C�*��St�����xJ��E����ƒ?H(�ɽ]�������a�?ؤl���䟝�,�Α^B�`w����ʶ�[�����kR2 ��]�a��ɡR�΁0��Ƥ�ʌ��T`xB�K:��%�R�.Z	K��T�P��%�x&��j|}�8�kSf����eЌ7�6���#�@�0��P9��}��ʯ������]�ף�A�,�Vy&d�z����m�x�(&!;J����	FX��K�>'rE~ځ�Oy�5��:FԼcS�����?�D�J7i�8ߣ�|ߖ�+��cN��nF��1�|I����EUMf�IL���幪Ƿ����F��B�I�KV<u�.��̒�^O�G�:�3[��٣�}�o�"�_{D%S�<�T��5~|�Kb�u��[�JLc���B"e�~ʁ���R&��QZvl�lC���n�$d���1_��:?Anxϊ��Q��D=V��^_�z<	:uL4����sW��ww���
Q�����+f)qu�@q2}ػ���u0"�Ou�>�@��^$���A{D�b�m��a�h2��?�ȻԣԾ�$�~#j6X����X�v��1�{׆���7Wl��5���MX�sO����P�7[�yȄ܋$���;_�2�8dA���q[^f�aƆ���.�������G��@���=�d�V��#�C+8�o��~ ��#Ѿ�c�oP�{5}dU9w�^��_��2/�����Hϴ�1��c[���Fw�IOG�:QGy��_8�;z�:eqӲӪ_�6\m&}Ρ�&���k��=�'t1�e��5�amĥ�(�s/���9�#<b�>�o<�".�^�``����9�����%��X��eP�-�,JՋh�F?�D|�'���Kū�4+˭�I�L��O����l�=����M�P~O��uF�Ԙ�[e����a���!��32_�c��R/a�֘�,�hάa���?�κ�1ǅLA�~t�L���IRu��^�58�1r+f��|���P˰���*��W!���/oŞ�:`���o����	�J�"����U&�G{�,�y��͞*��!$N;>_�54�>�'_/�O$��zc4"�PL���(�PaB*�K�s-�L��:w������p˂n2'�%��6��I���������6*?3��{}X�Ȏ1�II�p�G��=�h����_��O�}n���D|n)S����~)�q]�������$zlI�.����#o�Q���C=��h�eQ6�'��$��:�� �)$�L����q��#��o 
*&��s�9�e��ʴ�v")3�~i1�u�о���0����'O��PȖ�wf��3��e�a�0ɞ���VX�1�0�LX�1�0�)x��xs�&0�d�E�0Üʎ�?����c�)��i�9��9.`���A{g�:
��h�Ӓ1��i����iG��.0su3���M��,j�a,�h 1>^�������c��`Q�0Ü����cC4��'�Q���03����a�9#H�K�=6:E��aÄ�:��B�� jv��9�Z��Z���0�@_�Kս;DO���E�L!<�>l�߃c��6aL���Ҋ�o�}�2szX�1�0�L�U���-���F�&�`��P`����g���z�1�o�� �1�P8���J�<���F��\
�a��F�Ye[�7�S6���������=2(�}S��� {��U����1�+�_�l�L%".�H�$M�#>?��,?*^��2��΄�Z3��LJ��[�BH��C\^@�oF��j�/Ϸ�^�o���&E�2�Fl1c\cm9���$	3јLF�㬪���Y���{Ҡ��GE茅�?h�z���0#�ä��"�w� ��EȎ9���譒�F�!?&5u䍊/�#c��9�wHU'��+[�%YؙѲ�wgt>A(�-���+���L�?x��.:�i�V�ۣs�L��h����P�x�S�ʛ�a&���|\y�"��w��ā���d�C�&c�1Y��B�L�����:bA�l���Q�l�O+Y�
�4�-�"em����qX��;���r2����'���%8R�y�"OW�l�|�}��N�&kT-ϒhͻ�gzP��'�>Lt�v�OI��m���b�aƏ�B?r/�`O���,@��>�w���[T-W&���]�Uº�h����6Ǉ��4l����A7Qg�/F�^E�D�O�>�囶�C+ZwY'4�h!_sɳ�H5�1��6� ����h�!�8�a�9	�#���^�fD�'OVbq@:m�&���%&��$Ef���Kb6�ď��Vt�<5uuΌ �Wz���HCO�$B��7��ƸC^��n�#���S���+�׏���a�����ya��k!�W��5o�'$ގ�劮�(aK��$��+�����]+��跿a�:r���J�R�3nr��������|�3��םy��|�=ѳ��D�/^��1���]pguC�M�`f�P]נ����7�"�#�a��8�&�^ז(ۣu�q]�M9K��
�p�zد;ۧ$���$Ywt��D�g���0A��f���ѵ�#tK�(Z5��!�38�&7�<��|����C褵]��+�k�c��g���|F	��*���6�a�u��kB@�ɴ-��4��s{[;�F�0c�?��d&���5�8����-H�Oս�2QgZ��y�G�:��\�&m�y�x'l��t2�F���uD���fQG���'N�A�:�n�/��N�J���֢��&膠X�i7xa���	)�*,簿���b˖����ֱW����T���%�����?p:��k�EߥӯFӎ�Q���֍��r�g���e���he(�0�OBq`B���0��A����IV*ax'|�T2��z�>k�ڥXM��j��r��y3ЍU�J:�:"�L@±��\�ё�@��%׸q�'�a�Q���K0ZF��M����|w[Z�ꎽ����03Z,��=�g�,t�����%GD���F��ި�/�M)���vD#¢�<s$��Q6*-�}��� FND���Vz��F��"&3���귨/��L}(kڑ0�g��1&~��3јL&8���~� ���"�)ʒ1)�=}���w��2QrM�8T��J�s�h�}�V��(�\I�H�>t���j�υ�~�O�.�F轠�}!C9%�'���MG[1��!�$ٹ�03)))�Õw\�z��X|8k�W�E#9�%�T��֗zS�tz���#��umՄ,U^μ ��B�?�b,�2�hKl�e
�#&.�RI�7��_�^�#.>i���K������]�hk���3���4�K<�{M��N$Fr�|�C��4Èџ
��z��+qr�:�a��Ж2l]�����T�
����ȟ��������K��/t�?|�o8�aű���A��>�熟񛐘���<�ѷd ���QZ�� I�k��ϽXB���,�Q"F������4��jTz�T���,ն�<C�ժ^��eK!�y�O�ۗ���P��Vw�q�ln�􇌵V��+�'��|�W�n�8ǗD�h�@^5*PL}�>@Z�k4�0}�B�5�"$��rL(DC�Q�۵�5�4�yMc�|��2,�0�V��{���cǫ�F��@���/W�-�چ��?=_��}^?���"��k��`6[1��Ř=g��O9&��� ��|͍��8�,с��W˲/�4'bRC�3:��=���aĆBu根�o��!s!��k���g,�b��>�2lsj ��(I0���3�P�.m5����z����0=���jm��'��5�K�֭NX}W�s�_I��{$�2)�*e�B˰�:��K���C����K���ə��#�]n�Le��>��o?	��O��R���V�aqj����}���Ǎ?��t_�7�yDK�_ڼVٹ�pъ[���0M((��lGw`˻OC�_/�	���[=�%f�����o[�>�]�Z��'{�Hol��gW�?��.3�[�Y��]�u�z���:߇��&���ޫZ�;�Q���#���?U?�2��5;�Н�fu��_v��֗^�/�ǎ�uyw���n*6��KW<m.�⋊�N��³p�-��u@WG�о�4?lI>x��,z�w��x���c��%����$�N�0zPU[����;�O�aO�O��/aO-Ѧ��S�g"M\��l�Ys�b�%�U"�L?WY�}��ߣ��"$�
�4H����~�e��Y_��-k��皦)"�����u���,��SL�.DH����P�ԮS/�4x�!}�[�7��u�W�V(8mM�O��dx`qً��f��]jl��<ˏ���/I&k�aK���+�$?�h�1��Xy����3�� ��5�:�8E���me� ��
���6�ӵ��+�-�|~U���<��:��v��{rN"
��AbfZ*�P��V�'��7P�� ��M��	�Z!�P��L�y�^z���ػ��߅u�=����h ��C�6m�����۶ׂ�Ͷ�uUU|�޹QYS���/�87�>���L�e/r�I3�h�NU���9�eR��<t�CA�����j�6�k̓�o����7x�D�M���UԑR� MH�]r�5�!��x\v�W���_)1w�_?׃��b������":ns�a��P�ێ��c�,6��}��k�`4�>�m����{�6>�7J�z�?��Go|G�/�}0ǈŘS����nA����Rq�����{�b�fQG1y�%�\�&�o����}MT�!��զ{��{ײ��*)�ޘT���)�R�ي�d�cM�Ca�"z�����{om?dٔ:[��ݖT�W�t]��JX��Ӱ��)���Y��g-¡����P>����Y�g��f���)٭'r�C7�2	">5�z�Kx�_Ɔ�|p����{㱍[�ud��H,��F������³PX2�{T�C�Tc.(����<q�Q��J������aœ��|�v5��f����"ɚ�IKٿ�(�~�J��d�y�(�������U�W%��������}φ�Y��Ԯ��8R�T�Nz�D����ӓy�]��>P���H�E�0�*ʷU�}��1�Zo��*��ґ+����G7a���^k�SaO�)i�ɛ��9�?�J!QG� �����m���h6=�x����Y�=����@u���C	�� Z&���R<ԖD��C��'�#��o\ͦ�D�p��ֺ_���uπ�L���45��O-	ڲ��a�DH��ȼ�g��-�������~�=�zD޾y�����/��>}���%M$%g���j!;�Eԉ�ߎ�fa�So��jM�������ؒ��H�%�]��z��nqo��8�қ�uF�,�T���X�l��e��b�͛.&��Xԝ����[鋳a���EGW7f�q8��(U�����@Wx��O�x�(JU�_j^����x�W��m�k�Q����'�81�U���aQ'
���)���T�h�C{�#�|Av�K9K�M�GI�U��(�N��e({����6��U�����s7�Qyj�1jlk�/i�ztZIN�Nulfj����z<�	c����L\�E���m¬��>��N�~�u	�_�������ǯ��羡�ʍ�����{�j��'�#$�d	��b)O$��b�|=�uau�o����=*w�:P�d��;���t]��t��t�>���3Y�/2}�đ6{d
���d�Ξ��0�H|Zܰ��Ӧ�S-�����/���ߪv�ჵ;���t9?�u��v��a�Gf�WT��2�b�]U"F�+�^�Y'��ӄ!��^Bb9��qHx�������"%Mǃa�QI|Z��˷W�?���s��aeNhIv��R$g�P�3$fWDm�б���Hé��0��"�7d#��B�$ŇϛϠ���<{fgHߠ�O0ّ!2> i��~y?��nW�R�No\b�a���<�1�LE�/,�{��f<��u���kU?��?V��{e��cߨ�ؚo>��������{P0L��z��>�ʙ���%f�>q���l��DȈD �ݐ$2>��$���{ ��=�L	�~#��$�1��V�})�$�P��߭�"<b����!"���Ml;�aQw�����?��4�8)i ����9I�VT�m�z���.%5$e&���x9�M��HI������l�D������3���c��[�_��8���W����(|(hP��Ѫ��繫�Q)k�7��ȯ�9H@t$��jf��gR��.~���u��z�f8S}BQ��$u�.#�8�Eso�y����	����T��[�E���2~�k)-��+��7����ģ��ї?:&��[��q�o_�g�~��?z~'v�q@YZ�;+[f��NC\���.��z�|�2,�K�鵿U�m�[}����̰���UW'��E}W���^��I�y����.낤�힥��F�閸\��>���$��7G��r�?>�����?���>��y��ړ����&r<�$�_qt.Xr-�f�fO������ROt�)a��,,�E׾��&<^l{y���M�D�����oďW���Ǘ)��؋?#�����dQ�~��Cc��WȂU������p�5�rwi��b���ҷ���Dݗ
�'���$ت��+e�D]�	��o�e�	!�l����nZS�����B����+�-��M�.r�	�ϗ�س	�νz��W!�<_o�~�r* �J�NBoX]f��d�|�w��w=��Th>NlR��_oǚo?���V腧Պ�"�k�}=�ۊ�/����{t�ǯ	��ͧ�E����ob���TGj��7�6ܻtM�#[&6��{����,�ZzuwM"Q�WoR��"	�9�$�T�������W��L�	��v��8�~p�FM}���D����[_Ga�<$$�_#���v��Ho�EsbH4 ������΃}�S�IL�p��;1�1��Ș6vW_��t�n�:&������iG�,���=-nt�-��E���v���&������-dMK�}/|�z`>|n�.��n/����u�͟�K���=��#MjL��GyK�N�����w��X�/5+���-�>WzБ,�p��Ú�>�K�p�U\�zaEEKV���u��3��/}����'��������[y�T׊��L�R$%JP{������$����������9���:l��/���k�˲�h�*�O6/5�
G�˿5W�x.>�D�Y�X~��{W���'B���q	�X}�W�}�F{}':���ҫ:����K?�,��|>��ۍ���@�K�y��M�vY`K[=z��?a��w�lѾ��X�Q��2������|{���-�A��敭������֒�yG�=g%�_�Z(	�|Wyd��iA��t��:�ܢ�>�V��}�j�}ׯ�y�C��~���e��Һ��R�hFr�t�"S�ZQGtw6c���U�܉�8�lhj	��+��'،C�<}�0�0�AE�Ͼd���C�y��v��(ٰ�Uh��@w�Xl�W�uDks5^}�w��S�aw�B���}���_����߀�0D�
v2#�B�P�'Ӯ�V�b�vg���>^����;�.y����+��PDZ쮘���[I��Xb˙��Ϲ3j7Z߿�x���O����t�W�~��l2�$���צ%֓.��?��Ȯrr��ƈͷ�����gXt�gP:�\��y��Kؽ�M����|�}u6�8��d�Ӳ��A�!tw� '3w��f];�1��d6�dA��i��҉�9�0	.P�4U�����KnBA�U�H�;>Z����4���b�a3�a�lk�gA�y>�nVD\���0PR��}ϝ�������i;N|����&G�gY��+�戉�c�z��P�]W-�(�m��K���B�J��u��Km{�_�+ួ�>�+��5�RB0�d�K(�N��U�������'��F�Nr��Γ���7���;���ː/��Α��ȳWY���n.�x"�'��nz�,��*?S��������Ԏ��ו*�����i��㻡��@�@q����ώ��rk9&:P�����P�t�~���߁�n���dda��K�W8���:�Qyt'���G�r���4o����8hF�\q�e�a��ns��ֽ�o3����n�[Yo���B0�`�d�O*�����ܷ�tB��JP���6#u�k���L���A������y{��R)-�:C09���v��ݦOJ�^�����DT��=������d�Ƨ�h0*�{�[�.���i7�2�C�`m��dZ�hH�ƨ��>�S��N/��o��'%�+Ň&Z(��Aۺ�)�H��V��f_�+�`��!!=y���=]��ii�iC�,	f��kD^;�(&�lQ\\�R���}z�Z��j���l��G��=rΤ��+��Z��	�f���"Yk,�z���$k0{RP��;����
ꍐ��va��l(^�A�,ZJ�x�����6u[�S�4�ڍ6�^�����T6=!�i�f+,ёI�03�	���Y��5�m�3��Uw]6���z�?�M�kw*H��1�]�>	�TP_�{V\^�	P*{B��PBe���_K�Y�{Q�e�d�AI���!����xfr���(3+Iɳ��?G�ڍV��U�=�ft0#�(Z4���wm�o�E{�a�3Z����GX��w��y<�b��VԹz=x�*����x���)eܭݠ����8hABq �%�e��V�-�X��i�e��B����[vűmhJ٨�`�3����m�E���n��,Dk�D�����0L8�%?~�_�6_j	���͏+�����3ۑ��4��o,H<U�m��� �q�c[vX"�J�}Îٟw)M��Ə�譍��DM�����q�[8;4�ՙ�U�P���<ߛ]Q�A�z5&y�0L���
	:�ntC���q�u�/���$�{A����B'
� ���"g)i��vL��f���_��m�]�'�YZSq@���_�֜��T��%"��'�P��<�ϸ'�a�I���v����D&�	y��6��xH)��p���3���Ơ�|�y����^�:���X����f��P8wd$Z�}��#v�%�����%� .%u�w`��a�� �ᾫ�:o�3Z�΁�OO���6��U;B��T�����.Z�VO��p��v�&^[������ez�'���N���^�B�k�q����:0�τ̷��>@6%��aN�#ւe_��z<u�`Q�DYiX�B��K%�u�?�q��2K�p�w/�<�\�֑&�rW-zۆ�#Aw��o#9�x[��s�����2�������=�������{����"��ѵ$�ܚ+R�C�a3jތ���V��>kG�,d-��o�^3j7��|��"��ۀC�r��
���}D�ҝ�:��<����@�
/����������V4~h���af2�T֪�;���T��Kw�:J�=o�lT�������q�C7���J�M�Z�Q밅���pq��=r��J�p$�����c+��m�����p�IYo��"6{���2�[lh�59b�u�l�5���H��C�bI��/���Δe��8qA�T:��U;z������=���4*�)}����03y��mJy�!�=�W���Qq�lW�͌Kn[t���v��.��m:�7Z��C�TJ��b�S�B�p�	\�d�p�L\-�߈#kȺ@B����5�4�7h�w�����F����L=�R������N�J��[�׈oܱ͗=e&d-��*�נ��N������3j	Bp��]�)d!d
����hLt�TݻC�=�yjZ���i��ˋQ0g�V�^���#��f,*Q��FѼ�a�w6vCO�&6o���	�K$�h/t�ҡ�rZk���<��)����Œ�jf�QoЊ�RWDq�ܩ�]�����m�|����!Y��,���z"h?`Q�w���4���mP<itP���Y~XÙo�I�%G7��1��z�x���9�;J0�FUu�}y�{W/��������]�>��.�>�~�w"����!ȋE%@�>
"m�_��>X�Hd�o2�C������F������Kz#i�_s�r�4�жߌ�#�I�1�%)��-V4|`U־�x`ln ����sP1݁V��M�6+ˏ��~�������`��;Zv�k����7���2�0Y:껆��Q�����^=�o��Ms���eywHv�h���;�m��=+��mQ\����˳$
]�F�֙��V�Z~EO���ڔ�W��~y�A���e�:m�,�8_��7Z�J�j%6ى�j� �v)�Ę0*	b�7�5��L�~jX,߈��M/M�,�B>y褒/��4l�>����e���H��� F��.T��f��I1�Ġ�lB\j,z>s'{�"�l���`m5Z9�8�8W���Q-V�M��!�&����K+g��Ks%���5L�հ���SAK�z��f(>�6�a&�0�0YF�����Q=�o��U��V���#��0_t�ʸ@�G��:�a��H��v�+Am�Htŧŝv|ծ�a�=��\u����m�w�<|	X�1�hê{�9.d�~��k�ۛ> �L4E�yX��EP���jpds���K+HE;�c�S��h��ȇ#�Vz^���j<:��Xz��6a3,�f
a4`�Sߗ�n�\�F��b2	ݻf[x5�(��DQ���(�z���W�����P<_���zO����S�0��E�N(�M�R�S��0L�qr��d]��%H+�E��Q�抶a���D�h��T`�?>��S�����3�`0��I9�Y����0��E�� o�q�RP�����|�ϸ�7��p��"��u]��]����ecק�%]���x:����Y`�H���a��~���1��c<�R��?^Ct�ы��6U�����4R���߾/��ck����o|L)(�==Ce��)�ZO��^ϻfި�/�Z��~�nľKo9_96�Du3�HT�hsw�`����T���Փ_]�-�چ����%�c���C�v:��+eϞ̦'?B��T�E݁�I�8;����`�H���a�9#1[���c�)K�'�̝�x]y�e���g�*|NǪ[��d.g�Du�0�K��L���AF��јs�L����a�[ ��i�g��SXz��`�H¢�a�9�!����{.�a>ʶV��`#�孻��32PtN>���a�Ug'������˘0��:��BX�fL[�5渀�)1ݽ����3�ē����+�T�o)�A{M���@u�T֞;VY��'#wVrg�۬L�X\��~e��`\E�-!Gj �dj(���,!�����R��.#ڌ�'�T[BP�o��O(���L����>�U�'��( @�P�������`���ڲ�>|�V�}�ݽ�뵽�:H�dE+Y	$Ad&�<ӱ����{j"L���35��=OUuթ�����я�
���h�����{�-7��{�R���lܸ<n�@O�I 1�x,�����M-m$�GP����4�n}��vQ�*?��O�T|����k������%頡?������#yz�_��>���O�/G)�4|� �a�&3�4*2�+@��e��BZE��ȬR!o�YU�3�`
 �f	�JLO5�a�EV���T�^�I{��o|@d��`p�۰}�����G�M�� ��H�;:F� ��|��f�h�7W��
�	s����a��$���t���֡�P!�Ld���Y�G��f�ސG���'#-�Nt����E
6&0q�/d*�0%�& ���->$��p�'��3U(Z��d/>U`_%K��'���ε� �p&�O7|o�Y�	as<(EI�U�\�p�ݛ�0�"��@$���0�q�
�ߚ��hƫdy��"t��P���N�����)<S��dv��{�`I�o�C����y!���fo�B�/J7�]��;��6fo��!��{l��&�N�����04��+��%&˦��#ۏRz�10T��M�y
�<����rf�WZ_�A'����%	(Y�0Iv���J�x��m}�����mu�?V{]�`��ws�A�.7��遤2u��ho͵q�(M���I����uh
�)��*���['܎�N��������.q<��1��>2]�o���(��pC�[^H��P(Ҡ�Z���O(f|6][����wڬ��"�rf�P{�l����G3�4h|�7%��9�*T3{%��؛�P�`i����{�� b��o4F|9�D��S{�|�V�FP���٢s����|��|Tx���� LF ����s�,OB#�W�8��"eQ�k�x�a�m�(��OƠ��~#,<Y7�e�qsO&�D2�L�=�p	;� ^��K���.=�_0��И"4�c�w�
�0�Qv�l�O6(b1Jy�I��GRuxq�/�a��<�9���?���K�l/^���K�.��g�c7��9y�AĤ�bE�T�E�s?����&%��وN�,f���ǜ-�,�������9Ͼ%��B�qi2o�
�O}b.�;��qca!A|A0��`�]�&�"Čf����t�uQ�L��+mg���ѣ��l��*ܩt�`5���b���.�Zuz��B��LX�<�����`Z�	��p͕q���~�꙰��;?h��i�H�NF�n��r��c��g_zb��]W׬�����|x�˧_�l��Vq��T�������j��g�jPz����b��F����~N�[�a�p����IR����C��24�do�a�q�����[L�m����c� ǂ)G�uAp�"�X��P��7���8���j�T�	�&��t���ԥt�-U�

'��@����>V�\_�3�͛���>�LA1������� MpC��B����
O8�����q��8�.��\�C4*V���˥q�>��e����n*����n�gV�/N�^IrCi�l(,��`f.x�>��#���F��iI)�	+q�� A1s	�h�� ��M���菪!��������>�Ao
����8��C��\G����Rӓ�y?�wU".�5=.2��}�2ʓF��2��x�N�K����KԈ ][<8[�m5���Kq-������oU|��/IUI�\Ä���V���X
1�˟����ԣu؟�j���τ��^	s���?��� ������$5���ٳiu^��|b�2����n�d�@.e��U!No�:�Lݻ���p:Qr��<v(���j�=o�!�N��P/|�����&&��W�0(�U��Hc�ѫ�����֮�<���]q��ɿ}���Y�XY�&��'�y�K�/-R���S,i�oė��>�V>(r-��A&�Z_w�T��߯oyฬ���8���o����V�{U��Ok����[�m�E��6��!��u��E+>	^���̬<8�����3.�W_�5�wp/��(D�2�����Co�Ȅ�%��nO8�{�0sxsȬ��з���s�d���W|�9�F����W���Hcj�+�怽�xA�߷��o{�Nj�o�o|h�G�Yߵ6���e����z��X��_k���<��N�F��9�:Ӣ.�kQ��M����c@I|�g�?���g]��/!��,�Q�W�7�?�s�x��'�Pu�˺z��<+�}ѹWù��Ľ_n^	�r�]��s������di�/L@���uA3��zS��8�cb��s.�ޯ��
n������?���f�}���1�,�B���3,X��Z���1��K��__��Z3Q(}]��C\���G]�us�J�Qk�L��JN�t�aJ�����G�z�����_���*�}qY�����U�|\�\��O��蔔D�|��j��[t����U7~�}�_����k����:� ����!��_�-^v�%A7���ko��z�G02�˵o�:6X��ŎVr��7x���f]�߅&�}��a��K�\w�ixa�'bWpE�P�ՠk�4u��KF{]����=o��x/����\����~*��%�?���	��\��|����y���"IXqݗ�O�� �����`�}g��;��� ���7_��/zTRV��_�����[q����!$���!�&�D��c�UC��0�$B�V��5?���"��Ƭ5�����`���j��ŬZ��:ΓN�D��'���Gs%�;�����G1����{?׻M�Ur�bZ
c8��<�/r2+��ο�c ���R��.������`zџw��Q�5�#&�������)�ċ�Pbx41���^(��4�}xH����OUH7�b^��;�L�I���J���ػӼJ��k������!��3�^�Qt��C����[�������y���͘���=�S
 P�'�OM�K�庖�������Ƚ�����'y��0�N�9AN{�/��v�p�e���W@���X�DG���&��k�^lz{�(A8���R������e��/�O�UTσ��r[���W0Q�6��L�'%I#���m�$����_6?�6�Ŝw�gu����IG�d7����'~��A�߂�(����6񓘔hn�,��io���`7>_�+�Bk�n�����0�� ��2<�|"gV��a�U�j_�fI��6��Nbl��v�g�A�y>��x��F��N�u
#���w�F�+}o�;q&�L���X�|�K�<���C:�&�\�.H�� b&!e����t���Y\�ۂ��8�A����ޟ�>�6ӽτ�e�u�gL�2%�\������j!&1�Í��d�3��h�T�,���>� ;��}]T�J1cDݨ~5�(�!#3/-璓Wµ���u"���b(1���	~Ӳv��G��dc�I��C���{�d���	i@M�	1��s�����1<�+�xpI�xR ���P~w��	�JN���)��#;9��w�O�N�3���%��~�=^�
$>����`�e�Tt���4���-�t%��[�E�3�_'uI}�K���ą��H�&.��L\rC�G����-��H� 9��7�Ԃ����x�FU4PUZ�'�>`��wO'x�����]?nd�Tt�χ	�Q���L�7\*Vw�3��˯��XͫP���3�Ր���g{�by���?���6E�Ð��v	�yh
�:� ���������H�Ӳz��GE�%�� �H�K�
��L���9�����:5*��ь7P��[Y��������XU�r~��g5bM�(h/����mK�����+�����hMA�6��d����0��n5�M?�?B��
A]+�0���'�AY�;<��V֬^�/�q�S���N:>$�7�|�5�N������lB�$?�U���Y�ȸO�Kk�.����E���]\{(!�Qw���a�M5n��*�f��70�� ��j�
���O�6�}��й�JӪ�����fAd��å�Ι������_`~�6�NDz�W��>6��'39� ���RfJ��Ȯ1��ysTh���k�'B@����䔇��d�V�Zul?���Ɔm���ی�rv�ֲB��\�$�Iԝ�}"̹�����|�D�r������`��u#|�����`�y7�$ٗ��xp+�r�k���5�c���o_�@��������,�8Q��junޜ�Jg�F|`�{�!�T@��m���b7�@)Y�֨o��~�	�H~"qW�r���:�
�&�B�"�,3���$`��ἋS���`�����ۇ=T��RSMA�B��ٳ��X,�����^m��5M�Y��q�h�5�bz#o��U9�+[x��|er���7=���+C�^�R�+B��F��S�.��2D������$`����W����G�oX=��u�]Trn�_��|��H�h;+��\ƾ<��w�5�g��Sǃ���r탂Ϊ�A�3��x��:A01VU{�囏|����<��}\���%�1�P+���0�-���J��{�����;���u��^~a�Nw���V笒�:�dB��f	��̫g��7�����ie�=׮o��ޓ�Z�����V�/[�pʃ���Bq(/�7a�6�O2	�<�K���߂��z�chi� �l|�{�pkzz��5�A˶����nԀ�}@N ���w���[��h1����/2���
���z���oA �m���l����gC�.r�a��"������ଛ������J�����A�V�{]�"��gp��2�N3Q����u���{�����o����U��o0�߅����M�Y�Ϫ.�����p�y`��K�!�h�}�'pՍ_����c�߽6��G�T������[�C3�xX�7�g���a�V��#�CWO/�������H�)�%�}F�i揮�q%��rQ���
�����4����T���%�,n���xu�����V�����������5RO[������J�'�s����H�3���W~���{,�1�}"������׽�}=��ï��qr"�c�՞<���g�̲�u�	PUNm)r�}HF,�p�ht���O���W��K��{�c�� lz�Ihj�n�\G�F�;A1�5� �LH�e��~����_g,��#6#C����?A[�5�����hK�
��K�K��9j����F�;��>u���UU�;�ܰ�1x�8���tM ��M�r��K�fVXk�ܳ�mCy�}����{����
�� ����}@�g+�n�
�9��W5���޸�mQ����K"���V�L�	5
F����^�3�>�����MR�`��a��0{�2��;
��@��2�ca��<d9���}��(���7N� ��>अ�^(=?ƽ��&��O̙��kWPT��Q�����8t`+�4��^-GS�Nؖ���h_�v7�.�o�����R��W�v��,���w�+�
� �<Q��N.�.Ο��dc�4�1 -���C��+Fڷˍ���>p�_���
�2��E�	F����c�����Ĩ=Q+&@��l�;<N<1��r��3@�xA�E ����<���O�DpSJAČ���-��W�ƉFFa����� �$�=��@Q��5'�g��R�����*���l�Ea�r�e���*�N��v��1���[�f׶�5/��x̲�=�`��;�XV���}m=�a��U����2;���eJD��M�N��K�&��b�3q~����v>�F�6��ѻ��s�4MgN�!7'\�l{��nM}pF�0:g'��d�*�8��x��קn/��a���z#��2�*N�;�1�!B��n(Y�_!�V�g��ψ��I�[4�"��;
fo3��xJ QG&��۾�����|�ٗ����nf�U�5+/2��֧a��|���;#͒��Vx���/@�_�n����	�j%ȟ�b���`į��_'�ҍc�D��m/K�`5�0t�����T�t�灌rfo�sn,��-Ω�!� �O���59'J������Z_�B�8	�<gث��_�F�ΉX�;fFz�g,��6N};�н9}��)��\vN:�i`�d�23A1=�(QÓ~��ww�t��o=L��v�	��Dܘ1�tm�-W���3�e��O�`�mq��O݅�놶�ҿ���>�7��6l7��%h~љa_� "�`�aß}0�����	;@1��v�J�{c�'� �G]�:/��ä$7�B�, �7� �l�>!��O�g�M<惺��S��ܻ�	�7�$舓M��o�p;%3
���%N[Z�;Mݻ�D�SO���`��}��a�-q���>#V�)p�Lo�������X\�k�k�`��r���o��aO�I��Ū��W|0��C������&��Vf��~�|	g�Հ�WX%$�(A8YN��w��`�a��>(�0E�LN�+�Q��M"삽�@�e2X�e��6���69���C�{ �)B��rZ���Eh{���)�s�^��B{��Ԁ�NXƎOeA�a0Ǯ�/��IL�`�Y��rp�+�)���ڥ��!�*/MS��rv�IF�ή�{�����>��H�(�.Y�8���[�L�������l�Wۺ��q=�F�(:GA���Fv��h�E����]` ��<�0tP2f��,Q�pQ$�17�α�,�+�S����;%ț�B�2�5K˔��3gv�u3}\k7���ܹ*䣽�Ǝ`�F"��t�g!� f&�C0��o���)�7_�`�f4%�~�� ����+n�^�=�{��=lo���B�5xpLoD����X��@���6^�˪� ����xs����� ���E�tH���$���2g|Iho��hoA|9I}�ۋ0�!D���Lą����3��pέ�n�yP�q���{�AL5E����3sLoߺ�:�q<�G���<IȬf�2u��x,g"$S!�=�D	1!�;�5�)A{{w��.?gUbp����a��X{qiU	�ݨ7Ƅ��ֻ����=g����5^d���j���X�k&�ɫX��������a�3�^�9�}"̾����8Q�D�r�2���P_�D�	��``7���#��v����d��U���w����z���<l/F!g�����-�&����I@L�q{���^� +B�'����=�e�AA� H��BMhд�w���`z��� ��h8b��g�+
A�:��A��
l���	�3�WQ�a�9t����W&�w	�89$�� � f $�� � f $�� � f $�� � f $�� � f $�� � f $�� � f $�� � f �&�$���$���������uc.�O�\tA���nqZ���e����:x2�'�w���3��%� ����!�Lc�W��R����0_$@R@����?t��������uCoH�7<����1{`���_���~׌�iunv!��)�;G�@Q�]Љ�Ў��O�M���7J�k�x�Fʝ�B��|���p������KFAVpg$��E��oa�k�}�	���1�;�$M���dzc���E1��0��G��*3��|��iZڴ�:ov�)Px�b<	X�Ş"��T�����6^Z�ybg�ނ3UpI����eת�K�	г�}�=�v �IC`߄�"]��E�@������P�����!g�j��(�0����_�y�W�J���;W1H91���;W5^��[=пK2�K�[E.9����³�_�!��޷�	��w=��s��F�Y�D��e	p�h/���ޢs���>&��&��������@��BD?�<a�F-�K��?:S��^�'�� �+� �.����DT�<�Tf�=�o{���t¶�ͬԠ�8x2��i�M�;�^�����mTR��z}�u��+�.���͝��}�	�T{����	���o����t���Jk'�.<���i�=Aӟ�Z���)@�B
ꆏϛ+A���Ʀ.��Ě+eC��2hoN=���#W	O�-���\Jϗm�Ν��
�6Ƅ��Ȼ�l��&���OC�"�L���ƿ��<�TՇ��Wބ�J�!&DM��$I0�A�t#T��#a��QV�
�>�A�s~�tMn`5F�Ų��5Y��\P��C�x!���ԁ�D���.��ܹ��Hf�ʄ�>:8I�Qfo�%�{C��K���ޖ}0�z����MF0 �y�G~V:�{�ۮ���|���A��b�~/��Wױ�U\X >����C�#0
w���Rc9y�޾~���c���΂��#?�bq��?6��y�Ue��[Ww/$�c��ss ##x��P8�C�ǝWa~�#?���`xd��m�
����݆��a�݉(+-�t�;�`"��۔�m��f�ms��(�?�u�kg׬��ޓ
���d�8`��(֜�cL�ya�yr����^�\&�&OV����g�&�ă�O�
��[Ϟ*�?d��vS%`�A�T{혽$������K/<�s8�_���㶻��K��=*���������*c�u���C�0���O��E˗Bf�w���m�q��n�f�1"�_����c��7��=��#?�ut�����m<7�|�����x��0�0眵 �ϙu��}���7w^˗,���#?o߹�ڴ�m�_z�1B������[�D\y�ǈ�W����<f�kV\��Q����7Nue\q���"�78���3N=,]t�kF��k�/��֩s��ofB�i��[�1{�o���S�̺%��A�ù���'Qz��
�q��BG��!Ԟ�]�<1����殾f��T�b	� ���ZO���o�q8�x�跚.j��ZA7v�@!{�Q?��.��TXu�5*�,s��9F�ꮏÞ�@	۟X�9X������1���M�:��"��g(� ؁?pl���!{g�q�	*�W�� �Zȶ;6�����JHǽ���w��ޞ����C�=�fv�����x���}��������8X���c�;����������ݮ/�x/���}Y'�������w���K9��ߖ϶9�$���c�?�u?r.��fa�I��az��O=(�
W����ob���F;.��`J�©t�`c�M1Co`??��-��Xrm|Ғ2͂e�5Wǡ�I������^#;�˹k������@� �T�-���MHN���}t;S���mN�>'DN�^���s:�{&���;�1Ot���K0g���:~�S�)�'��d��ٖ��Z}�N�@�\!ág}`'8����T����Pu��/�k�p���KdCP8��*�h�}t���DZ��S����+mw�BA�F�e����D�J4�N��F{҂0pT�B���?�`�p`���	.��""�u|���cG��.E��q�d�7[��,OJxS`x�*X�<|H��t����y��������L(*��̬|p�DP��@Og#�4�9��1����3oz� ����C�����/����PPT���?Rq���)	�@��m��,ǋ��H�X�˨΍�
	5��e�b���鍼�
M�<=\>�
��=��IcŸDNN�
&Qv��UF[�_��hi��6�=�W.Y��ߙw��I~�`������J��ԡ��i�*�˭���/��s/�	*��É�nK��a��@�T8�g�������e���7�у4ډ b�R�Ժ�B�����|�	�i�l�ƅ�*	ػkl}�H�1�����0�;��2�2KS�=��艅:�_.�O%���ka�����5>��j����L�cL�V��d�a���Fa�LEIcy���:6z��}��A�o�ky�����c7[��z�����ɻ�e�!����k�(���h-���JTR��˯��ˮe�p�"Q�`��Aݜ���ˏ@K�N�#�/�A�P&���Z� f������#q�/��Xt�I��8�P?g)��⯡�� �R������F��ԩ���w�:�(�o����	��e�'l�������i|��������^#/�������u���!QT5��Ӈ���]���Z0�\��C�	pݪؽ�����,P��
6F̬RS�S��?J�MJ/��s0{�2��y��ꆯ���v�͵�HB�T�H��A�4���St\�W]���=�{�@0������K��ƃ۸���1T�A��z�Y�~��]<��Bm�߯o~�f��y���tͅ�~R{��u�%�@q҈�9�ŉ9���M��\����0�Ͻz]�?��C?�J���	��,Έ]޼D�.xYv�-�ݑ�2Qx�埄hdZ�vq�Y'QG1�$�q��.^�iK�n��_���G���x@�kU�a!&oO:�
b �	�/�oz��c�}�H��;��<s�5P�'�p�G�/8S�'X�c�xm���w��5���ݫ�,]��&���U�i�&��۱�b6��x����s��o��0�%P"�}uf/-�A���	�
к������S>6
��~{�{F��Y0m�����
�{�<.��~���AnA�a�̡�7���x�'cKM�U�d��)Q�YəK�7=QAS���+�;��h�T\�0]���pM>���(���K>v5����pβka���Y\�$xrU�S/!�:"���#?˱�j�}�ܞ�ߔ#=�/)u��}����ո�����J�m���6�������O��mf�N���$�9'$:��u��x�������uG/�tG����p�|ؖ��0�~����یs�N�e�j�8�apߛ���n�<���FN�nc\3��k6�g�z��_��Xݭ�?#3�\t9l����}��:x2uH��}b���N��x�#Qe-����Y{��{?po/>�|�@�X�+͗y1%�0r��h��~��ֵ<�6�������ue˕o�����"��|7F����N�-8�l|���ܛ���#&����񚈝i�p��ְ�:7t�:���5O�M׾!�u*P�m}j�姖�}�k"m�p����:���}�mv��v����d"��t�2^������g��u�!��d�ٗ�_�dҼ�%�D�?�Ϲ�s�Ո�Gz~���/��٢E�M���vIG��3u�}�|�n�.A�=�H"���h��,6�7o��ʗ���B��^���Y<Y��BA���z�,���?�i�E�䨆��Zk?����E]L�旵L�~�o
rxP'MQ�aT"ݮ^T�`#���?w�Ω�0�7�ZM�'��f,*��tPRV�%���7�P�F"#p��r9�R� �d`�4v7�8m��S�e��_�Ǔ��9��.q��Z�eUp���x)��ҙ�3����tFbS�N���~t%,��l�;�<�.2o���BHY9|�kfiZX�`l޼NW���.x� &��y?&I��r.Y�~Ί�8�Qc�	��Ə����]��1���&�Ψ ������&L�Xb����!�t��5t��z��T��n��!3R�[���28��(]mm-��5ANE�z��\���{o�BG1�}��n������AaZ�9e&�ė#�x�f���m�����<���\��R�0��T�r4MQ��@AU�d���W�A�����U�>Zk����G�����p�.]`�����^OmL�mL(����C���e%k ��P³���&rP�8�B����[v��>���#��)��:�5�������nB���¨Z^M��d%7T�ͬ�t�$f��ֱ5�yڦ�K",�/�|h�_�W��uw��q_����s��qӡP�J�Da�I����[�"�z����W�W�@ bZ�ܐw��7���i�����J/�?JD�+A�	�x�"1�+Ԗ}!�&�7-km˧�l�/��\�2 u�0%��C.c��Yr�T<གྷ��A�	�$|�D� YS�h���7_s�)�;���e�>�щ�A�:��i_��X!���"��	(�{�GԵ��vQ�HĹ*_���5� Pl�;<wVR�v�7���l�}.Xʧ7���D]��9���4g�
�﷿1k����a�(��������wTYl�ZϘh�r����lf�}����$5�t����y}����bΗ�>�v�s	θIy`���Ă|�:��/QA؉̾�����%�o�s/����m�p`�FPU���X�5����*�|��O+���N���ʬ{+�櫟�u�g�KS�.�!B)Ǜb�b����旄d?�)���ty�t:C��k9��w3&�l~�iXq��0!u˦����Zy`�*\QwC@�f@pz��|b� ۈ�x g��a	�"��w���/��-Ǘ�(l��2�>��7+�2����|�#{J�*��7�}���H�����
W�#��)�i�5��M�k�7_��F��U��m��<]be��;�/���m�7���-��E�E�d���̡�CM�YP7g1�ʻo=	��*�X�tk�	� �2��.`W	�����M��;�+�xt����!�[5Je�Bh�wsh��	n�5�~��ЫV�����WW]�����h�s�$�D��ipB�,X[sM\8�d�W+������=�Uu�?]�T��U�go7� �q�x�����|��c���*����7��� bf�L� ��`y��>�W���o�� ����7��45l��/���]j!��|N.�κ).�������͊��Zݽ߬�,���Z�^,C)�k7�Ϥ��%���;-�my���U�zI$��o3Cw�<��Lo�����o��/�TY����.��~Q�˦/<�3����B��%\�ba.�~�����2���� ��y��\�I�1x����|*kr틽W�~�1ؿ{#��K�����^�K�!R@����g5>�}qer�?�?~l��	mVι���r��r��ټ���m�D��Y�	�K�uA��o��]�q�)��:7z��2��!���7>���mWU�W�pGv�v�E�\�����)ζw��!X�w(�^}����Ͳn65���6����[:ס}>#�JA�<"�^H0�����(�^xz�Y��.������¿M����^K�ڷ=�T���n(� ��ePlE6���Է����=�Εի�\�lz��ۮ���(%?�U��SqQ,�Ͷv�=��IL�:<���<Pw#���8�L��Q�F�����{��QWc2�.?�r���b�*w���N�`�_�v{�vu��Y�X�(�} ���L(*����<��n�����^��l4�\��9����sA3l@��*WĬ��l���������=
�*�'In���쁮��v[>O%&@�ԗ"q�h�����Bc��R �Z=�$�|�Q�ٷ
�nHD\M�"��d�/W��(�K�&_�u������ӤR���c�&1�E��.vv��/� ��_�ҵ�Z��3�$��]c-짳Ǖ����+]t��5�7��A�X�y oA�{�h���A��+]tn��6٨w��H��X]8�3w��/<���17�,�oz�$�%u�k^����l���������u/d}N�9y�G���w�|\�^� �i�~��~*
N\�	w����Q+}����X̑����0t�y���k2�Ӫ¢i�!�⵽��<,@+����t���C���Ϩ�%� f>�t�����h��_�Yn#v2�
�k�J�M�����Qf���\�$3�>pCF�y�R�F�	��k}�gD��A�.7˒F�j'`����(\!� N��x �4	�u�I`��kT����w��Q�Cf�3��@J�_|�i6�Q,��_��AV��/(w��M�/�Z_�;�[ί��N��6��YəA�$��=�9�ǌ��T�����?Oh����;b(�Z{���˾��+�˟��C�������	;���=г5��m|�u7��
��M��lo� A1}��]L�̺9>u�Nt};��1���If�1������my�g��s2)�V�z��W�܍�S+NZ^ex��]`�^��T}E�k6�-�f�q�k�h'E�� Nw�� ��C�qȝ5��H��2�
`�����-dMr`Ee���F$m"�3D����ט}��.w��b�.cMg�N6F� �_�U�\皇k����Ϩ."� #v�oX�@����N���	�Ȏ��&&#b��
���^a2�p����ٷ�d'�$Ý"T^.�oyR�]�����,�����Fｴp�ގ�H&���IAL��Ի���c�7�*=˱���֩����belՊ�Q4���0�޵e,��i��N���DyD��?� �,���:�(7��n������>�Ԁ9����Qn�'��	�B� � N�Ɔ'��]���w����ո��n���N[��b}.��h �f�Lo`�b{�/�9��b.�~���,�4���`���q<����.(hp��	!�^\lB8��`I��-ġ�8�����*^�lM�:�^� �y`k�A2^d�6\9�4���(�}�s;�}@H0t��[��h0f�j)-*�++p胱�t%�Y�.�xaWh���.�?__^�h"ztcR�� �	�ȕ���H�h�O7a�v��װ7P�1{��^m�� ��^�r�PC�Nz
"� �/��x�+`������ՙ�M��QRŢ ��_y}�a��>��l�M2^��`�R�,g�h�lW)���4�q��L�;�:�7�����TLJ)�ţp���&�8�1Տ/ �V%� ����H���Qo`~?�NG����\� � bBH�AA� H�AA� H�AA� H��#�	���ZRnd��^���1�B7xJ�U��I6��� �	��#lG8�+;OrY� �ϕ�A�$H�AA� H�AA� H�AA� H�AA� H�AA� H�)��� �ǖ�� �,[�Mh(.&YI�.[ki��������ʕ� � &�Iu�B2*4�����K�;�[��:� �,@b��!"="��] �Xs�S��/LBf9ګ���O`���uA���v��;��<l�ɶ�BF^����g�?��`cj������=�,� w&ay�r ��r�[	�h����/?	�\�~�G�Ꮢ� I�|*3�+3�!��Dxz�_�����Z�l�M����a��*���w����"(���ODZE]Fi��' w��������l&�*
A1���>� r��_��*��VA������v�``����6n�逪j�o�>������L8�4���烑�ؼy3��b7AL	��3�\�<�G�TpyN�D����a��J�³��o�	����u;^��K�竐���'���=��j��c�F�Df/{1�D�m�H��ˮU�tY�Lԥ>Q��/C�y2;to���id�jPrn2�R����a���0���	������Q4M���������8��u�v�x��x-� �7��c�7P�����%��B��O��7�n筞1{��P����f/�&���wK��읎�J[E�7[���eȪ�9'�}p����л���xAS`���b��	ȶ�^\��c�����c��	g?9$�Ihll���*(((��u������AS.3V�������3�P �};��Q�U������J:��@�B��x�`�>���mu(��Vȧ{�
�5E�(Fx��yD��.�\[�O���֠�y/�;��|����E���R�騪j�P(ASF�
)P~�l���5�0h���b�S���`�
鴗�#\9�t*�����KY��MT}�y�'O�{2u�sG������TUǃ7Q�q�_8y���$��8��u/�}0��Z#W555�O�@���O(�t�
K�$�£�ڸ�,0-j��b���Ln����5�`q��OG��/>it~Ð��и�7�'N.(&���A
����gr��֡����C7٠��H(&xvm�{S�����x"p�R9A�ɫC�-�s���b���8�G^#Eh2���Y�� P�Z�P�̺)ͯ�``�����C�1U���90�Y~At��lI��1�A�용]\�p0�t����Aa?(��J�=	���d��vX�;�x��)�쭾2���lag��j��O���0X���]0�/}�\�'1�{*Jϓ!��OA��0qQw}lj݇��DyTH�Ҥ0%M��HB-��A�͙���YaeVf:��U�BG�iibT�,t�����sA�wz$oA�S�T����8��*V�52��]z�j��~�S��jw�{~�̆�ܢ�#�_� �a�����w~c9�.�w\��������k����]�@A�,�>j��G��W����G`g�N�(Y�<����5W������u�"N�_�A�"z�ڷ�_yi��_p"(���$`t�� ��1���:,� U�P��]��_���@�ڋ� ���dW O��`�� L7����G�]͉Q�	�0�r'��ɺ`�^�;W5�
Z��|��J��R��봔*]����L(,����<v����	�Fh<��{�,�t���$P� ��K�<�%֗�\�U5g@u�PPT	��\p	"(�#�=��y����04�e��%`p�I%u�[p�b.����I�9�x�� G�fAG\�ė��g�$KQo`�f��_"�;����u���#V��k��76�z�����~t�U���tm��ȪQﯼX���/�[�(���*��[7�8��� +�����x�Ȅ��z8{�U��~6����s۬������KA8AСxI���0w�rX��zC�}�G�@�V̆�ˮ���ݰ�'ax���H8Ӽ�,z�O�ӚP��b�[�o����$F�5���/�8Θ�����~����:����� N��œ����8'Zg�L2*TK��8N��%�>t@z(S�呞�#'�v]�C��|�{�/"�}����7��5/Eg�е�z
�89X�/*%��\������>��t�'���<l�+�1s��ad�Iաqj� �2�
<VD��+��"TV/0�Oe�B(��o���߽����{�yR�mϛ��;��Ը ��y�P����<ֲ�����-�c��+Ż�o������g���,�a`��CV�L�:+՟(�>��]���7?�����k��M��Vi��Sc��e(\2XdO�u��u,��(讽�N(-�Ž�����
~����'��u���A���&� f�uQ�}�� �p�7 ���{_Qt�%W||�����\�b�*�J��f��7��P���7*�n[����f�[����?>��Ľ[�(�?Eg�c1%Οu�OSW#r��.2���|z�[���&��ìk|��+�ժ'Ŷ"<�Z�UQ�%˹���t�^�YK��Ü�x�F�a�oq�Y'QGL+4��8��$��"��ԕd{
�T�<�ݵ��JH&�0�7 ���'ݶ��
��2m?�'	�R�T A���lI�}�e�d�#���#^VEF�2���/F>�SQ����!ӂ�������	��z��y{ҢޘV�.X��\?��C��0A�{H��ᾟeUi��2����| .�bkp��n�b�����-{at���>���!F�)l�M<t�6A2k�=C__�)gK��]�1����)�`�I�������G�@���K�*B~V�I�u{$���A7�^���^H
c_������N���% �Uc��|�h�Y�@y�\�.�E+>]����,Xj��q��N��v��^�lMЍ����?���h�g��M�YR��nL݃ܪ�m���+��6O&Wwmv��
9��>(ʂ�I�t�7C̨�+ZϽ�f�IrÒ�n��^���}Io~�}ΟK8�H� h�c���pʊO�T/�"x[s �g5Y�x{���������;���,�u=�����OD(�/:�A_D6ͼ�a��&l��P(e�F��d�h0�3f����v��Jx�3���n[W[^8�g0΁�.P�cBQ�4�J��UA�X�R��d�/�ҹ�^X��zێ�˸�ν6��'������C|�?�;���b���-ҁ�j�O�R&v�ٻ�}M��	ӡ,���#N��jL�:!_�K|!��7���;�������o�K�g��� ��U�g@fV�	F�6��Ģ柎�9*�:�4:��`�XQ����Q0����.�U�9���7��O^8g����{'0�}��?��<tJQw��+v��p(*���de�~N?%�Hb6�a&���K=����>{��,86��ю�,��C��K^��-�t��/k�Xk�L�φ�ۿ��w����|�L#Q���e�����>6����FZ�5y��n��`_��5�g��`�V!س��>�,�%�A�q�W7�0�\�`7�L��U:����3*b[�v��Ǘg����7� *n��؈�~����5D�1�S�)Q��,<D{���?86�M��޻���A.��JI��_&���X8��p�:1@	u���e$�����z�0���Ȅu��)UU�LN�E>��ҁK�8+�9�}���1�#��A~�iS<��C�7����U�qJ+=oD�e��:�_8V�M�:��c�0�T� ����aZԉkO
.Έ��K��dd�=�ak�0�s��?92�K�I-	���:��$�B�\~uqf��z1E��>�R�ɯ���B���4���y�E����t���x�,�H��K��s&�?���X��R�h��6�K��x�]#쯦�%�3�k�Ňi�� \i)Qc~e�g{��R$���m+=}�L��_ a�S�I}�n�G�n���5��XL=<	�n�,�?�uIL_N5�?�?�>X���Υ̿���?ӢNH��fB�c�4����w��`�"-��<�kR�0҈s��G�tP�Hn��E�ڞ&JA�t��t^����	���,�-���rb���nzU�cޭ��ei�`Li0�7G�����g�d��EF1��Pݣ#}�WPv3:�ǵ�Sn*� "u�H�.�^����hd�l���V��ι���1��v��o�=�:Wi6�$'`J�%B�9D]F�V����,�ϖ�o�XU{����@Y�ȉ���ɴ�]�iuݝ�\۫���4Fq:��N��@
��G=]MP;k������W�(���_�`�9���0["X���2�����������k��c\$B�H�Ň\\�cr�п��)�W�D��?�۵Y�&r�ab����M���3/;�%ݶ��\�$F��Ϝ ��*�n.Q�#��u�/�[�Y��c�e��ۛ;GF������;؄�X������5>4�=�S* �+B�,(�|��7Vj��W;���,�����Y��z�~��o��� }�)���0�v�Ý� 9$S� ���Đ�ģ�C; ��L�*�w�xè��u��og��u�s�|�������QRdU�}g,�oxoL�D�����s�,���$O�~�~������~Q�T�R,jT�����j����sH7�?�p�7�{h�	��°m�\�$.㗟 ��9D{<�����ɤ��ѓp��c��Q ����>���rd�M����W9
��]�(Q^��e?�)�r�Jw@�Yp6_�

Q-6��_#="�q$����j
�Q?�J�����z�+g����W�o�)�@FZE�-v��H�0{��ߠ�� �x�8{�U�
8�1��n��AA�b}��O������&��༔���4x��_s�CF���w��%l_.��L�F��o��۾��G����i��%.�x�h�s��ͅvؽ4�_�R�H��2F�\%�X���Z��~ª�{WW_�X����})D�����s����x�@̙���a��{��?Bk3_.j�A1���&�6?d�F�������π��3,�k/��(��%��ƙHj� ����I�5q����+�l&�~ʳ�K�H}����.��@����9�O����n7�������o�g�*�A�o�ky�y����~�,�����J���Z��CuG[R[��g�.R�g]},��?�s�]g�o5����/��k�8j��.3�t���( ˲����K-!A|��&~Q�˰�<����[��s.�i)��ꋿ�����F�S�\��u�;�֘������V/5�~����������̾-~n���W���g��!�=h��e�y+P�>*;?�Эo{n�SZ�+M��j8�c|3\ˆ���EO����/=_%���Ӟ�_L���ǄavoE����4�s/�	*k0��L����ݛ`��X,d�\w�AON���p8]]]���1����� A�u{�� P�珰���p9���o�Ҋ٧���ݹ���"$1�B�f��ԧq�%#'ޗ�'�p�A�
;�����ӫ\����xI�g�ZX{�;P���䫅 ������.U�c6���o����"]�z����A�����[q�>$���(ʷ/������,� cY\ʩ�,͌'�o�=�P��j�+Z7�@���/�yy�ugÐ�I%�gd��(�Ȝ,�=�},���iӆ��>CН�H$����*�ζ��&A�t�g�jo�0��z�=�ĿAN^	T�,���*��\"oq��1��T
,��g��e��=�]gm�tf�s?���]�i���$���+�b����˨H��5ZJ3�c�"58ku��l���[�7�ڍ�x��P��H��O����6:���6Y!��2���X�7v��� ���:������"��(tw�:"���mmmF���vN�A�T1�,�H�ٵ����`��Jm�{@�_�<!�$�!Bf%
�8����P0�f_�1)���'�UA�ᖘ�oz!�J3��y2�����fM�+�go�]4D�M�(�n"6��PRRAĘhʨPAt��pØ�C4��y��qU�N�{$�������� M/z�����k�>��*ϴ?g�z��b[�W0�4c:I�H 1$������җ$��	I6��{7`w���{�~��!۲��f���s��K�x���9_y���%�E�!+�s�{,��-{ځY��~D
O��}x����3�ЍE�b��h�oV>���+��w�	/�~�^�	կ�Qtqd��CAի��81�X�YaA�vr��].R��ēxz2%��m�!��9^?P��C_��%�Ql�G�3����!�d4�)�j��V�����9�V|�e��9d,~�9�|N������S�}������"s���`��}�3v}�_85���o��I�E���T<��n�@�<9�;�p�]���7R(=?��{;�L��]�C!	�	�(�{%���gOnБ�O8���T��x�����=�q-�:[#�C%�P''0U/��P5YAG���8&l�I��v�9'�I~�*�@�~$�V�������γΫ�F\nK�AzM-6�v���4T�\{~[��u��Pg�G�ĦI`O����o �g�ijB�����Ԡ��+���{��υ�y���<2b���	�`Ў��I;�/�J''��\
N<�@O]dw��+��;��Mj�M�3}��S}����W����)�C��k�d�6���@'��.//uuu�;i���	W�����3,E��rS��ՉX�xO2s3��1ǧ[mX� ��ƶ5�)�J�L��G���å���Vx&�SS���'���0q��L�ҧ��5�+2�Qz$��#��nPHB��6�֛Qr����g�=�?�9tgӸ���	[R���dh��i���222�p8�ZuR�d�����������&���ˡ�}�	����~ded�z�D�`����yq�v�jmD������2�^�<IG�D� ++�&]����U���k�늎�7d�>�c���㑽܍i��0�!�ʞp���h�k���0���⑳���	�u�mh�gY�H!᭴�T�&lp��	�Z����̌b�sg�Y�9��V��;��DK�?U��4�74Ci�I���T�t�n �ʧ�b����>S���ߙ�ŋYK<a5���[�����]uA�\u�X��څ쥞����B��7lh=]mRH_����o��M{��\�I}9#� ׼�QiYV����"g�;��+�3r�7d��ì�#+7٩i�獍�c�V���j�E@GboN�/B���kG��D /�?�R:�T�6��{�"�>��=�&8�+�N����~��r>������X"��c��/��T����w,��6P.I1���Qokn5ia2��ӍB�F��j�kC�
-�-Mؑ�N�{ڣP����}ڧ-� mNh¬L'k�m�w�R#c��!a��2�,o��M���W�������+-�YAG�!nOB��5��$+���x�7s}�~��E�'��v����D�TТ5�-��c��7����=e�+��� �^�ф�����l����[^0�u��-V���y�xh����i�٩p8�cFa;m��SAՋv��!]o�<�6�F�#Y  d˯�
sD��>�R;��+����6[;�,c�+�K�V���(k���m���]L6I�>}�{�
[�_����U=����c�	�6����	�Qv2%=l2T*���  FdIDAT9��|/�.G�_/�b��v��E S?^z�17�JDD�C�Kw[���=K�����=��_����Z{�8���IRP��>��J�m�@n�)+,r�>8���ӎג�hM���c�c��}�������b)�'[�t�cJ��F���Y""�I#�x:˴�(Wk�D:X:�G�\�P��GM!��6���î�-�T5FN}Fq�����"y� �,�:�yE�;q���!!N��e��9��׻�.s����h�1�Ѹ��Hv���An,iiiX�r%�|� �o�c�����³f������RSMAA�,Y��SC���&C��CJ=���ē�n���`������h21�Ѹ��.��za�Ts��ڱh�"��f�l6C�5��`�J�,_/g��'&$�}��!#-8�s��Œ�DD��h\f8bNl��*H_o,�	o�mύ^j4�;� 6�hy��k�U��|R�3��:?:��^s+���&CQ`�#"""�uDDDD1��.x�>D��j��80>�N^�����A����s�7��_�s�&�د��(4���#Om�B�ɪ¬=�ɦ��R��a��[�h�j�h�l��Jp�K$�;�G*����������U5��:UC�=.x��~���B����5E"�v�hm�I�s�sk�MBgF=o�1km���ycBB�5я��>$���=M��>�'�ݣ��nBo�	=��Ԙዌ�b�5AE�v��>�e��H����x��M讶�����xp!""�-ُd�-J��=��_�L9���x���)�Q�Yk��K��QǞ�^��׎U���ZG8����m���z�����o�B�IK�鳽H����� �+[��]|�7+<z��8aF˻V��,�)��K��A�<�^}����9ǣ�����U;ޮ��>^""�L�+���E��H�={���϶$�=J�!�Їi+�w�t���oO]d�Gr����W�	9g��H?�d�x���-�!w�GA�8�����U�C����nL�B�%a|������z��������,��.�*K;�l�x%���Ѧ��ꗾ&���Y�i�DDtv�ff/�����#	J����֬�GV}D)��k�Y���K=#��!���=�E�����#	�wH~��N�SC?8�0͏����PgA��v��&��Tz�
/r������l�x�u��b�x]���DD�RfxQx�[n5m�}���,�~�O���d���b�n}zW�%M�bv�퇭�~�o_����	u���v#O� �ǞR��|�ͮz���#�t�0�Ǜ\���|�|ю�Ñu�4o��/����5�/fӫ=P���l�����foP���}�n~"�p��N�k�z]�����7���q|r�#�*�Х����y��&}�IZ\�]���k7���̼��y��I�k�N�eYQ��}B�yH�k���&�t��\�D|�5�YC$�R�9��:���G]	��x�DD�$S�f]ׯ��L��0�*'��P��x���%�1�N82&�x�q�{��~��m�=���q�:k�v��G\�����[����X�l�����d������5��r�1������&�<����L|c �Xy��J�/OLǊLs��ז8	yC;��j�Fv�:�IZ�3��
t��{ԯe���+N(Y^��uY>�d��:Q��#b
�đޣ��;'%Н.k�G�`�y��$�g���irV���B樓T��:-��$���Ȩ�'c��N��6�+@ �v��8'��{,s�pu�#����BO�Е�dZd�GYK<�o3�y_x�_�~4��aY ��5n}�f����x���s�a"I�y.�hq8�ɢ�v^�E��標�IDD�'À�ّ�M_���pI�jE�'t] 
����lF��>��P'an�
7"��}�/s���B�EB���"�x���}��[�QLK)�yF�*�̅��Ca��70�y�+��%�7�q���:��^�
M���+Z S`���+Z�K��s׸V�������� ��W��񯶔I��\�jx�3��R�/M Ek̥=�Xlpj��3�Ǖ�`��	ՊX��^�.4�+)�NEߵ��aۆC���,sG܊XC�.c�q���7U��j/7u�7�_�]9T�EQ�eK�ϊ��K��O���d0��7�i�5$ŉ3�3����O;�̚�E3!+�P��t����ʎ�A��=���{��д�
Wg�uQh�NM��5X��ɘ�`
�"3{:��S�__jO���]�,{Gk��{�H���5$�z�-X],�[]���4��5�_T�j���U��G�~B�m�l�=��t�ʹ�}�H-<�)or0�;��m�w[�v;�MJf�[�n֧z��M����lo��-8ߵ(���n��l����^������d6c���X��RX�#�	|E3뗕�]��[���`^�UT>��:"�X$�tӂ,.,�	��\�K.Ђ��Cb�f�Z�_:;��֫������0)�U�u|���e-5���~U��]n���)��Qq|��xxX����M�\��g��~��$�ڳR�6{�7l�4�p�K���,A�9�����h��@���x����,��	���Ǝ;o�^l�E�E.��-��ֽa�7�Vr�/��E��q�5��S�}��p��"��M���C����pɜ�Z���9gDDR�*��ԓR2���H���>)�ٸ��;��K��ƣP���\��+3����G��z`2��&y#��ف�o)���n��~s��ᯛ�6=r��ק�v~7w�GQ�l�A��i���u����������ÎVg�z�����4pWuK��~u����N�s%������$F��`eq�q�I��C_�~)��zι΃Ñ������o�i���i_�-Qh�%%g�Z�=�OH	�,>��	x�?�Hb�0�2Ç����m�1�x/��#sT����~U~��@�����d�|���}^����unC��$l���Y�(zץ+T^��Iʞpx�;�����n#���+��m���+i��y�������Y��5t-Y]z�mA�A�3e8�j��1C��͍ꈈb��+K0���bņkn2Н2g�t���vFH{l�����K��݊������H�;�/+���F�n�KW�Zd,D˞�Q����.4���-н�q�R���Mw�[Z��#Ŏr}z�]0]�������,X���f"�s)ʏ�EsSU�������[�MDDA��^F�����А�XV�{*��AWGs��I.xo�AC�I���ռa����_���.�aK������_��x?'�4�T(�@�1�=�P��o��JRs�N�q5��������?����R�U΀J%�%L��xz6:a�b�a���_q��x��_~�@�G�e""��ۣ��$,\zQȞ_V�._u^~���ǡ">ӧ�5*�`�pw����e��w?�P{�k�i���BOB��� ([��:'^{@�..�X�n;j��_�і�[B�o$(�p�u��G��Hz���	uF�W�(]��f��������ր���PGDK���5o�>�J%��������/��82T-���cy��E�{}!Z�p_�=�O�kK�Z�W�Գsd��P�<�P	�8Ҍ�)���U��GB���HW��^��5P��g�~�%z
�/����|��@DD�C:'�G{$�u�������T��h�K5�7:��}.��y����1}Ev�T\���L��B�5�؃�7�ʶT}�!�@�wk���k��^�`	�p��pa�r�,��k�g�#"�2���0�w]AFVAX^��sFB�%���bS��|��������<�-�N���{v~��+^-��j��p9�V��o�l�խT �}h��Pgr+��]?S	Ii�no��y�DDF������ay-��#	hF��{�L���j����Uڴ�ف��!���5ԙ$����׾�Z^�E��J�����'-*�WR��3	�ӷq	蕘�SGD+�6-&S��Tm��KQ���0٭JQÓ74�z��٩��%������lQ�&�?��,|A�j&ųU�%�3$n�S;;�C��\��n�n7""�@^���	�ۥ� ax[� m��A,��<^�7PQCS����Fn)����R��d`\ߞ�-݄M����A�M�6Y��.C߼`C���tw�7�,��m4t{�>QlP�����iɢ��M��jm�n�&�>�m�9N�%�?!vKѦTGjW���DJ�J@��ա�2�@!�|5��Ľ�x!R_�^7{���dwgp��R�Ɩ������a	uu5�����PGDK���#-��Wڣp�:y\#�A�Gbe{QC���y�_����O D��Z��j��1�X�k7�|�>ۃ�=��k��,��S}�I�n�M�o�Mvj�K4�-ˉ���}�B��߃��Æ��jc�:"�X"�#-����͞�:��Av�hn|�#�l�=r��TI��E�1�ǴO7#D����FK�8ۣ(��6��>/�M��#)���o��Uw�8}����o������U_���Y��[��� v��C�|`�+����������""�А��)3�}M�a���"#3tS���~Fj��������#9�$8�3�R��)ߺ���w��4��Eߺ(ki�#��!���h
u������]�C�~�q���[v����7�	��,�z�d5�-;���mq��[�=���M�+�F��قw��@Y���m��CEDD��������7_yW_���,��N���2tg�Yv�
��zj�6tE��A�^�N8���^�˛1��%�P�)ٞ�����ƶ*�m0��O%g�i`�Yr�ݑ��~L_�^W�j�ϴ/���)�~篊/w��̕��E:�-�`O	�x�[��`w�E7b<�^7^|�7�Gc9��b�'!"�В��u*��7ԝ���Oa������.W^z����Ev�����$#5�����Yn��v�����w�y^Y��������܅F��x�7�Jҕ�v؂i��-��^�0�o�])	׭?��I�k�o)��H�w�v�UΛdOS�Z�/�i��]c�x��vG<V�{MP������S��ό�����k?bA�c'��w<�=��]���>��<v:;�o��:��HJ��� c����_���/6߮ܕ?����ͯn��Mz�����Vz��[������DN��+iyׂ�n��$���7U�l]���[_�Ry��g���%�\�����+\�q�ƫ�H�b�����"w�F���}�9tu����o����j�m�����R�durwm�)Q贼k5�Ķ���������a���AsS��u�z�Mz<�7��:i�/q!.ÿ��u������<۽n/�����ޟ_�ʵ%��6�#��"�P'ÑZz��&F�k�I.�-��i{�s�w����(��9��Y���?sI����*4��\��|<{�gE�BO��޶齋�!˱�l#c������j�b���3�\�li����]m8��%|g+�~�=���m�8fQ$�k2�C|F6�t�����<�e+.ì���wRsu߮�q����̬��SO�=ufCU(���a�����wX�|A����5�/�%8�>�ٽ1wS�)�=C;�+�y?����d�`�6숐���c�ϰ~��� ޒ�b�:
ֺ�j�vmo��n���k�{O�=UER�q�~�gn�,hQW�|�$����$���?���O ���9EHLJ����������'�[&|"�^��C���KDD�'�orqP�cow;���Wl������&&��b����чX�]ks͸^co�	]!�_V������C���w*���Z�X/+j3z}�
��4;z�d0��'�z�z�����&�F���~-05��I8X���r�q�GH�תz9t�VRw�i��V_*Z*|�hgIr	��W�PC�oE"Y0�vЂ��G�ɼ���%���ڣ��R�B�֥�
�xM6U/y�:S�R�p��𣏕�K'w�Խi��MC+C'J뻖�ʯ�Ez�RK�:8�429���^�������H*��qa�H�OoCh���W�z�:#+'J�+�["��NN�2��I���%��Gzժ_1��X@�w�M}z/c��9��/��E)mR�����z�y8�7�P�F�{�<=
*�u`��P"��N���m���7��"�6%P�wE�-?�'��X8���P�ŗ;#�x��9�wG��!"�	#�Bz�d�z$���p�q�=�=�"uoِ^�ӠBI:TN<��ŉA�=��������}��H��:���$C��
.���=���.'"��ԴG�_?rW��'#@>��cZ��2ʪ�쥓{��>�x�oo�v��k@�q��O��\A��/ن�ģq����иۦ��L��5)]��C'��S�@GD4�սa��5!w�䌘I�:ɚ5�ڵ���br����I�T��d�%&g�n%����&E~�N<7�op�~+<ZJ/Ҏ�b��㕞�O:��+��[�����m�5^R���	���OYU[�ծ�
���D��!ﲧz��B2����M(��i�Օ	�|c[߱��5�v��I�q�?�P��e�8�Q�����{��Qt�-1���u".+�U�|V�^������ұ"�lK.w��lfP���R�?d�9�k��_㐹ȋ�s]0ǅ��RG*MO69ޣ��[��u��CM�KW�l��"�Ǯ}_=�8�N����G�����q=���ws�6�U/)�	�DDAj��s<r�����sF�d����z;<��5z0�˵�]�	K/���1Q�ˡ�"��ڲ߂�Cfd-�h?`^Xǟ�eΜ���2K�
���ٓ�����]�-�+g]r��',uv�r� y�V�:����f4w�!��0��_Pz��_ѕ�� �͂��M)����V�'v�YK����N���6}j$��Bi'�X��ԃl-s��3I����^�.�5o'JX*��
��]64��e���Bo�������Uaַ���yd2,*s��b�����������������3g����2¬ܔ����}����b�@{��Kք �#�@ݹ���Hj�F2_���<i�m�J�H��E�o|�yC:�����E��fa-�+?]�f��aOQ������7�T��?�RsM&|�P��%ߨ���ptU���������Þ�M��2� �U=y�.�x]���/���5爈(DT��L.���>�=���dL>i�\푴��M&���6�s'���"�r����#U�%����&��jm���x�Z��@�������G��S���Ԟ��I�ў���(�I-Wg{m�F��W�iJV���a"""��PG4��(X�9亲���G�������S��=N/��5���Y��H�9�p��Չ���c�����y��όU9PN� ^�}�#/��9,��$k�u��󌼨)1Á�Ҵ�_{�>T�i�ug&#5�Ա���P�m����KG|�}#�k��V�3��K���d9u������љꈦ�T-p]��C�{�Okam事�gᢍ�O~��Ћ��򨏿��",������ߪ�3?;���\Rx��co���{G�φ//������ww�j���+1�1�X��G�y�2p�����Wi����Q_��uXv͌�_K |����~��Q��T����c��GF����_���AO�hNl�љ�Ȁ�N&���WFUU��U���h�I�77���0+�˙�J���!��(=�}0�bg�U�q��""""�Z����QԲ ���hK� (�������eˮ-���7n@kڝ��|E�.DDDDU�կ���c9_�I|�����_W�E�!%Ml�Q��a�&l�U}��*�ʿi�n����(��X�n36�Q�ǵO�8�����^�p*#"""�������m�>l�lɷ�����*7i��
"f�U�Q�4�..ɆĴ�!�]��K����MXZn�v�S�mm�����>~��4���'���2Q�}Ƙ�)w��Y���'s��&g�������F�U#o�e��;�+�r!��l������ku$��<֜����N~]�4I����f!>�q�녗ڵ�(��i��C�	;����}�+z�z��}o���/�%�+�{����}�b��U��K����a���o��m��Z��2��%"�(Fd'j���n[�&F,\?'��k�����(�B���%j��Of�2v��������(Do��껲��~�tӏ�^�T�P�D~�Qz�ן�ܥ}������K�sޤ*�]
�]DDDDQ.�P7�მ�ڇ?l¦V��*ւ����&̸Cݠ�W�~v�]�}~�K
��h_�ADDDDa�Pw��Nܳ��������*��(@����(,��m9��ڇ/�1�k�������mȈ���B.��n��e?j�>����o����y��
� """����P7�7�h�݄M?�E������˄��A܆����(�&%ԝnp�O}{����*Tܬ�I]DDDD�$b�ӯ*��W���ۋ��(�W �6���YEL��@��*�_�8���P����(�T�<Ѩ".��R��N�ý_(���no��P�-@	|�q"""�)$bCݠ����mC�P���
�;�c����h��u��[1���|��^��OZ�� ����H5�n�Oj~�����>��wӂ�4��t�1�Xr烀�u�����
""""B4�:?���р�uDDDDtCQ`�#"""�uDDDD1������(0�� �:"""��PG�>��
E	O����wG���>7�����:
��-<�v�����6,6�H�������(0�ŀ�ummm)n��q�����_S���1+y�^�#"��e��ꗩ�����3�mzć:��y���3����k�~d?���+ ""�E�}t9�}j���+��W����PGDDDDg�PG3�MHHHV���񀈈��ń�UYA�7ez(|�"H�9�p��������5�r �HII��s/���r}]M-z�����/� W�o\�w���?6�DD�d�����Ҡ�
��b��`M�[����3�ơ���>mȁ���1>}����]� ""��ꈈ��b CQ`�#"""�uDDDD1������(0�Ű��D��&�e���O�����(|�bX\��ݰb�_j�40��CQ`�#"""�uDDDD1������(0�� �:"""��PGDDDꦠ���Gh�h�?���7a�5K@DDDэ�n
RUDDD[ꈈ��b CQ`�#"""�uDDDD1������b������}��p���׾����p$"5#V����n�k�jCsekH3�(DDD�KESC*��BKs%|^ψ�2�LHI����%((Z�}mF����n ���������M����OFJjń���=�_B����ADD�I��[k�Jjuu4b��O��Fz��[k����a���ț>�hJ�:U����(������>�ȩ]�a3��P4s9�r�!?�������꾞^����ͭ�7O~�͠�{�� �Sy���pp�ZX����ك�����X��J�/�L�P��T����F_O�Yo����'���,YqRҦ��5vV����5 """�ʎ���xUW����9������`B�'�˄�(<|��̹s��T��
N٦n�tݾ���1o�E(��
��+"N�+Q8����/�����ݨ��@W�>�I�v��$�� ]n�o__}ei��9g�E0��^풊	r���T���;҅����q�h����r�W""�j2�j�ۏ�8g��ύ��8����a���`=R��p�ڙ��J��G�}�����h�ï�����P]ׁ�^���$':PX�����oh��HN�Fִ ""����X���a���{��3������]�x����z�|L��|>/���b��u�_S�����ɯ��O��� �b6�I��{GWo���S{sKϰ�۹��)Xw�L$&�9ʬ��O�����%�DD��3?��/��H��[~�c;�A����Ј׿��b�@7����-����z'ϙ�L����huY}k�.KF1�j*߁��v}k{�]�����[߉G�>��_�	�!�'��!�`<�����L�V{d6K&��TA����R�͕�����DSKϰa���}�U4����ߞ��9<����ub�@7��ύ7߮��u���_]�A�:""�!�sgr�����-���uk�n�u�<�~��	�t1�z���svi�u4�Ump�}�ن��4nODDD���H@O��v?�a��j�Y��꒓î��V6[�AL�:UO�Ç^{{�>�>�qT�}.�?�zف����"CbRZ���\'s�f����#g�UBd�' 3}xo\BRz�Ԫ��P'[~Y��a�n��<��1�}l����e/@_g��y��\E����,��tղB44v���c��,�hm����/@���P'�3�B��KM�Cvf�>2%��z�홒��{����{E���h�M�y-lq�I{~g�����Y����:��\/a�����8V�2b;)cr��3��2|�U�-(^�h��N6�=3ԉ�$.+[϶XB*M���x�ǎ�%����sì�X�u�r-G�����|�muȟ=�K
P�t:J��!""�|k>x����0=��d���+���/�v؞�z/���X��UU5��*Wկ��-
�6��o�_G\"�Ĕ���E8zp+<�C�����B���	}ː�����r&">19��+�<�.v=����Tт}�J\r��Cn#g6���9<s�+C��=܀���?�࣫q�w�V߇�h������A,�p��7��vU����<���';�O|[�R��t�5ػ�1}�Ꙓ���pn��b�X�]�kǥ�u�Re�����!gJ}/�I����DW�&�Q"ɡ����R����\��ًv���x��/��3B��|o�m��^��v����&s��?D����^>�m�7�������ᄝb���)ڿ}������1�sB����B�
�$fC�((^�ΎF��1��K����z��%#3���O��l����z�����]���;+��m�n;�x�?�`֪��J�WcY3~󕇴�9������)$��L�V���7��˝>)�xg�3hn(3tߤ�L,<�rddE產�ub��K`�Xq��#N����-Xr)�KW ��7�9�:��l�B,�|�*�W��֐��?���G���ϯϳ����50��ڟ�1�Q��=;ۇ����;X)�AM�.wV6���ASW|B*V��&tI����ްξ�ok�ڑ�]��%K��;��;w��u�͑=ۤ��]O+Nx6��yX��J}�>V<��k�$�A7��ո�ֵ�n'���+��=�����ޤ:!ìsϛ��}�x�#�u2��b_5��L�Q��<����`O]Ό,�����J�\�����k�J=[�#��$�w.Z�Н�u�+u݆�h�?����z�B�w��v�q��S����h�����b�?O��Y|���:P���S�}ν~9���n�W��?oG����w^>�PGDA�qN!���O~�����!Mu4Y�(�X6eB��ɏ9y������l����ի����������*ζ��!�Sn�׫F��]�C�� 8�C<��9�����%�ePKu{@�N
������D��&�nЧ�$g%!�4L_��}J5{���e������h8�<d��Lf�YE�X|�<,۰ �K���"Ӕ��6�LH���T�\uj�Z�,�Y�>�mOur�٫G_$�3�ԙ�԰#"�H�U����ߦ�N�s���T��Ң��b�j,o���7��]�@��>=���-�a���������o(�L�P7U��֋�]�1���顮dI,��\2�Oui��u��h"5W�
u#:�Vہ������[Wb�gއ�F�H��_����	w��_a��߇�}%(r0�M1��j���X�/���M��3�8�h��=����=MM���:����o_��.��$��P=���g�E�?xsΝ�Sg�������C�����z��xBj�v��w���T}vwK7Z�0\�n�h�_w�m6�����{}�g/E��)Fz��5Lz�C���|�PWw��~{�ř "�H��X~�"����w]1d�D������o���[%É2���ތ���_����6���9>��"uZr��!��}7���1x���'�}�ݰəѳ�V,c��b��N����}r��᫁�y���ϥt�X�<E͡�C]��&��w*��ܸ隓e��߭�TR�����2l��o]ax���z��J����Q_t��B�}W|�"��c��bҦ����~`O�gq۽7����|��ɯg,+D\�c�ǔ=�n;U��=uD��֑`���u���T ����{�kǵzUz��\��]�d�1E��)F1)�T;K{�/�_���>}e뇾}%�S���?��wz7������l������:$��U���(�d8��q`^�C�4X �L�w���߶������v���`)���4��~���`�d�]�uSІ���͇v��a`����[ۥO��i�r[Y�p�_]-=x��#�0ƻ���z]�/#)=DD��H#�����K������oW����\���L�S7���[_ 1�z}����%�A���n
�����_�/mܳU�`�t⚯�Gb�А&K��ߓ1�0}�<M������!�O���.����BF���gN~�`�lL��O�#�@wh�1���x�||��ϥ1E��)j�����O���_qt{����aڛ7_�>�:�Ǔ����X� "�H2������L������߹����Þ����<��N��_��5�*djʹ�l}���͗���~zS�E����U�y�ݓ_�0�E��),-7_��gP����J0��$�K��
dޅ,����b��uz$"��S���=Ҡ�:���v2���wp�b���;��w_X�\����3��k��s�\0[�M7yO��U�~��{�N^����ҕ%��0�~�i	by�s���,�>�|�R�̯`n�^x��(\L�S'��1FdU���x���E����C��48� '�Sͪ�b�����ײ�����/���엛��=�����w�v�g;��g��b#��uaJ$�)G��-C��� "��y�����n+po���p՗.�{�*Z��"�&���T^�%Cԟ��Mx����ƝN��G�'=	r�����IdS��T���2�6W���nw�~?l�x8�H�,@FV��φ��S�ꈈ(�H���Si1D $����ႏ����^_4P��)�~�>�FܑKEM��8�ݝ�#�����/]�M�<�vG�KW`���0��3E�U�k��RK��hk�A<�7�����R��Y�̜b�k�]�Lr�&����y[>�g���] "��$�������J�;�]�+Z�rUrq�8��'�s�~�BrjN��bv�ꒈ�t��`��'��pF���8r�U�T��e��Ejz�͔	u��ZU���v��g�B�}�N��v�U}G���l̜��E��N�T�xt/�xx�^�I&�J!�t�Ll������ͰI����eh�j�w�p;=zͧ��^}
�$"���a�U��K�����[��	}=��G��mx����#3��dJ�:����:ڌ��']�r?I�KV^G\�T w�{�/��_<4�z	i2!V���|b?�|����c?~O��%�p}�.,�H�S���k�,>|Ç1�έCۏ����;ht����\n/:����U$&ش�ȫ~}>/���0�^r���-b>�uu4j��?����1�˱�����uEBbb�?��@w&�y�-î��%x�_���׃�<�g=ĝ�������~|Y����a�'�d��噔�=��ˣ��U�v`�;5hl�9���HIv`Ѽ\̟=mX���<ػ�1�駢fEL�:I�o��'-�;G������>G )��(K�}]z8�`�m�ڢo���d�W��֐�d����fm��B��@����CJ��m��Y��Kbz<��c#���{�o�p��
D"�?5Z�^x����ԧX�d��*�=P;��I����娨jÆ��j��4��eĮ����G4��P�b��gFt��[��P=ZZ%�\')}Zv2�i�fz��U=�Csp��Pl4�:�{�Z��,��?��!��x���3���ӝs�B\��5�yN�>���(T�=D���<0�n���M��!�����������b?C�dkn��W��I��_�z'F8뒟���.��x~.�,/�+��s� )9��؎S��t�8�t��/@�������'��������nKDD4��[Gn{���GO4c���H8c�����0R�l��.�7��;�T��δ�`=�X8wڰ��тݼ�#Zɒ�A�V���οqŐPwɧ�2�Qđ��39]^t��~��k��ǒ��!����Z#�Ŭ�����\��8\�c�y���<)���.T0/w���d�:�$z{'��(v)��SK�ͣ�a>��G��uR����v}k{|>���w��ǉ䤡�|�3�h�u��1%;y��%g%�:.)��R��h�OHի]��f3#+3�-=��lBN���e����������NV��݂)4R�l�):{ �:�9s�5����(����N�5ݠ�ef�TϴzY!�|� � �s�Y���`�rJ-b6��ǧ�W�����,�x|Dr�}�q�c�.�����]~�B���^4x���)���Yx�2x�#���m[� �����K� Z�d�Zj?3�I��K
���ʀc��{�2�l�""�X&�cg/�@vg*-�DNV�� ���C�V%�v
��'Ňs�F�1*'oVTmL��׬Y�����oz�T��v��yy�wz��ݺQ�cM&k�@7�(c���d��ŋ@DDD��d�*47�@K����f�vU�v|~?T?�>�#>��_�hL8ۍ	���Tﴌ|�N����[aI���s�PT����:�6t���8�y)X� �i�#>�٫8�JDDad��ʵƎ�Eksը�3���L����[�Q����dG��TY4��w����#�bv�U,\v:Z�F\�:-;I���?w���\Y)3����{����"��b��n���o���7��~��[�%+�W�9�<|0�'�VU�qK��V"�b:���	8�WD_o��;�ې���5���[oَ���|��u���"���_��r�M���B�f&"��I'�%.�����WQ0�̘=�}�͟��G��#v~��H�
��W�.Z�VBA\|2ο�ؿ���;��h.� �5�uj2JS���3��OU���1|�m|4�ɟ��@0��.K��^�}���0Q�3f٪k�`ɥhi�@[s5��:�v��!O��IFH�(�W&$�!��|��[q��h�;�����k?EAN^)f�Y����Iy�(:�q�Z �PGDD�$�M��_bݔu�di�\z����X���j8���r��Z��R��Y�̜�]a��mNDDD�kJ��A	I����t9��o>|<./��b����F�za��*� |Ń�&uS]|J��b]��&�f�������:��ז\��Ǜ@�ꈈ(&u����}\�\j�M�6��eNM�h�PGDDDꈈ��b C]��m�, <���D4��c�n�vK�++��C]k�h�gK�"":;��3CE1�:"""��PGDDDꈈ��b CQ`�#"""�uDDDD1������(0�� �:"""��PGDDDꈈ��b CQ`�#"""�uDDDD1������(0�EW���=A�W�� ""
7�Ӈ]�>�}��m����C]��݂��DD4~�j�d7ov6�;��J�>��Z��o��~P�0�QLRa,�%e$�u��!�=�]�ye�{jo@�=� ""�XU���jLj�����P����w���ϼ~c�]7*
b*���gF,��S�_(<">�#'m�J��WTtwu!/�`��w~�U����~�L&�CzI*�Ά����b��)�.�R��޳ܾ� �fuDDDD1������(0�� �:"""��PGDD�&.�ѬB�S���ƅ����&�#��	�c��pݧ �@��XL�p��-f(�r��P�8�*{i|ꈈhRm��ܧ}����;=Z �Q(ݕ�f$e&�d9�T/p�U���z\ :�:""��Ku���uZ�+E���î�v�����1�QD�}�f�Ƣ�~���c�#"��aQ�O���PGDD���hMz�L�quDD1�þ�q��8�:"""��PGDDDꈈ��b CQ`�#"""�uDDDD1 jC��(>�Q4P��~��u�ٳG�E��'""�)D�����6m9�����Y��M% """�`����sDm�өʋZ��4����"����SDu�SM��)��PGDDDM�+/��9�:�m)����K�ܫ�UKADDD�T����q;��<Qꄪ*��(�����"���z36���4Q����I�wݩ �@DDDITt����D<Uԇ��nvo,��SP����DDDDC�t_���'♢>ԉ-�l������/�h2YT���fWUUѰ�<�[�*�&��N�D�N��N��%&. �$�8��'{p��Q`l6۴ÇN��AC���:����x�7Q�3�������m�ή8_����h�-��Y�"2F��}�c�=�u���񽫤�t�Z*�V3LWl9����|ޘ	uBv�N��V��(X�	�5'�� /�(Z���SO=��W^Y��j��u)���vj_���*�><��S�N���u��ڹ�q�_jnQ�ɰ뒏ΒF	&�	>�}�:Q,J�z�2{����}�����.�}�t2MƓ�\�6��W���K�zS��߅�$���:Rm�{T�9l�����Ȉ���ʶ�691���'��؋w���>���Z�;DQ@�i���~�잧&�u�d��@�=?�u�7�n1��U{�o��@8@B��S�]5�v ~f�������b2�|���������W�����[ֿ��_��k�ﵓ�@�� �U}Jz��T����U�+�C���X���7���&�c�I��_U��V7D�p����Ã���;���Q@�@W-SRR�Ng��R����ߺ{�Ѯ����o��UI�dRe��	�Z�z�����D�lḊ�A[���E� �b~~��M�����~��D��C�) 2hͿ,�D\�}�����ӎ�̦��8��_;@D�N��_��������W���/Ԯ�Z�a�������6��m ���2��t�����{"�{�K�������o�l�kS�v�w�ʕ����s�ίi�;�v�y����)ðO=��+�D�)��Ckh�}>�o�w2(����s�ϫ��߯�� "CV�X�#-�UiA�=�ń>���5 ��0��54?�>�����L&�b�X�_�ti�((Z�{x׮]G�~�����o���JO��aX�Y1� î���&�#�V�A-���/h��"��˗�߹s�����_���uj�k)2��㏿|�5�Ԃ���PG��zȦ}�7�R�54����gժU�̊+Z8p����w-�}佫��]�"��Ó,΃ѐ    IEND�B`�PK
     ���Zv'ON��  ��  /   images/0755f9ac-cddf-41fa-8c34-4d71983a54be.png�PNG

   IHDR  v  �   �;ߎ    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   PLTEGpL������������������M��9w�X�����k��<�P��'g�&r�(`y'Ztd�2q�c�c�]�b�]�[�T�������j��,cw%a�h�m�i�q����&q�R�#~�%d�\{RpEf(Wx,Y6��t�)Ii"@[<a�Bo�Wz�Z��O~ItAv�1o�������]�����9�����x�ԥ�������������r�����������=p��׻��J�C|Q�T�(I;Z6R==5677== 8* 
!"!$889������sst..2,./MMN������FFG/E&"$%%())bccSUW444++,������������>?@fhk���������"!$##"000\\]zz{������������---////--! ������+.-,.*)3&!!!#8:) mmo���&*>Tl���009HXfo�p�����99R\o/0���Sg�#AB%"""���-+���*
#1 )8Ey0Q��6	�ꛡۇ5Q0";#V����qT�?&A ��d�MD�f���~r�Y3h!/B**K %<!��v,C&T��4M1��r2K.0I,@(C%/F)=Q=�ŷA��j��O<5*53VT96{��+uq64	ebIGb��4��C�Ƈ��V����n��zuq}�?:1��;:A��9�e^�qoM_2$�TIoC60��H0!5f��������婵���򘩿aNF�G�<�g   QtRNS 
#7^Lg*I��Ĥ���م�������]��������z���������������������Ζ��������������������}�o�   bKGD�a&�   tIME�7���r   orNTϢw�  � IDATx���	xTי��&���mǖ��%A:�$68v�$�LOw��V!��V�U]�V(t�TWK!�\mU���$K��J�H �bQI�B�c����%�ӝt������{k��I��h���~�=������o�e�e�e�9�����������wP��XD^�X��/��� ċ�q/���������Bǃ��,Z��/������{zP?��Ï<��c����ַ����&|���{�����D��b8��G8�ڏ>�8�}
F�,���a������O�5�1<�o�'�W �������
�{�}����������2�o��!O?�̒g�,Y�/K�
^�a��3O/~f�bB��o*��Y�P���2�t��Ͼ� _X������_=���}��;D~��3���g��O�?���_�BEA��'�꩗BB�������=�����<M�
o/�˲eAA���<
D������Z���w�"��y�2'���ă���Md)�N@��_c�k�oX�~�ڍk7�]�v�u˗��XA��7,&O,888$8xq�U���{�9"s@�8�JH�K!O� �g�<�>Y�B�+赛7o���#�g����7�]�| ���p<��z�SO���$����>��4��<䅠��+W�_��rV�����Q��V��0���aT*�� �GF�����q��U+CC�~�=���@�I����t}�>��w������p�0�F �j�*�F���t:��a�����i5V_�hcTz�� `�?��B�	{�� �% y��']^Zd7Ԩ�DSeX��P�G]k� �J�C�8��������h���^%+����']b:@��O>@�����@�!sB|IpH��A�BCW��)p4U�*�H7&�e���q��	�II�D&9>~���8����8���!�hxH��T�OGQ�_�|����l�P�
��gГ��'{f��,KC� R	_�~��qu�:\�Ũ�XF��BbjZb�)�O2����Y�$1v{vff�̌��$C�Y��X�"24yl�����7�E�/C�O�؆��7h���, wAsY"c�8|���(�Z��ł�9AL���Ĵ�n2������Ҋv�X |�A��̩f�o�l��e08MH�>�剄H'|����?��Jl��N�N�%!!�A����o���P���ecy���d�JK�O�5m;�=17��[����Y�5>��ؒ?QiN��vU�M��*�����F���Q�@s��U/��~���4��g៚�W̜���KIA%�p`�;w@��+����dT&&&	�5@]�5W�d�%j7�[�+�69�R�*��`L�L�� �I�!H��T�>�`�h�:2�F��\������	",���*y�<�0q�%K1�[	%x��H�y�J�� 4.�(
�M�yib%�D�\�fc�(�dl-��2$V�w�q�<����F4��i�=	~����
���W�� ��&����Υ��nx�����W`Z���1�������C���_wY���d
eE�A�N�p�J���Ă40�$kb�Պؓ�J#P�����i9%�=1�زE�[wd�	�&�`l8*mU�A*5o7Z�R��M�b,� z6�ձj�v�����Y?�3������З!�%KB��At��#ařO����U��J_�*c'���W�q�i�{����,C�(��I�ak����E� �&�@���*%�D�j��0-�l�ῄI�J���?����t*��pv�O-��g���w_
���B�
dÙ���[���v!-��\*c�$�n�lL��O˰d$��3�Ub8�v�$�$�WH��D��fr�A������E!��RZF����>�|�/�/(��E�y������1H�RQP:͉T�9�������P�ȫ~Y�l����vQ���V�������3�K
�NkR��*��|[4YMi�Iuu)j�go�n7�z�{��맃����yݍA�пK�/Y�8(,���B����՘yS)�N�K�`��V2Yy�����d�%������,..�_�`G��TV�:Q�.��bjZ�����ǠI�ott�޷^~yūA/�=��'�_�?���#�cE����!t�E�
��&�o~�`��R�lU8�y��2	��&�]�&A��-&� 6S�c)�d�d%&�v�C��*+��
?��(SǨߘj�L�`F��\���X@p���dv]����%�H�}��ti�x��L���\4�
����I0ƙ	u���X!�N�+���T^2�i���%ȗ,����	f��RГ�����_eM�^*��'%
L|�$��db,a�V��_^��_���C5�?�ܣߥe�{ЊuX �Rku�9�J��U�R�LL�'���tR3@���D���(�0�r�o�M'�O4�m|�g��\6F�YlL�����+±B��c�����?���B���+�^�$^�K��"D�Z*%�,#;��R��`x�uL����s��� I��D�$�O�X�y��W���B����5��_�q:.�����ӈQ���r�B�X)P�t��8g�V�To)�'2& 	ѹ ͆] %	��wC���&�*������u1�o���ČKq&]��H�����#����	sŮ���\�Yc�8�a��l�11��t��>L�����L����S��[o��-{�����U�����ah��O����@gr�RA�k�M~j�����
�N���[��0�f��$�I�'}�R`ֵ	vV�ըb ����ˡᯆa��#��G��a ��7��,ń4t����:��U8�X
��$�'`�q�س�*������l5���ђ�0Y08 �jXU��U�W�z���8y+���,&����X֍� SV����oN��n�TPR�h6���;��3w�v��A�)AL�Z�SGG�}y���~!���@��G��%R�IW�Ǻ.����R-uQ��]�.՛����b��(/�()ɨ��7vh �1I6 o�0��J�N�V9�zy%������Y���`^��cO|��J�UX��8F�W�+>t��$;��-�K�d�hw�c�Gr�� 3�m`��T"Y��(	�ʪ�i�&1M�SO@���KB����|�/KC����Tʲ1�����<��C�h+�����A�vC?�e�3���3X<�y9�����F����_B�������L}���|��䙐�p�I#�Ʌզ�H�X_,��U�\J��sR���\Vn�Э?�)v4�fr�Z�bmR�D�"!m}���OӐ�O�vz�(���.F0O�T��r*�N�5m��"ة�)v����czdC�H�˃��;���Ӭ**J�aP�Uk����Z��_/^�B�����NC]�:�K�2HJ#Ռ.F���L6cQ�Q�}����&v/:�-�����Pf�R��q��hW���\���W��?��i�K�/	!Qc�4+$%&��f��H*c������n���`j��2BpgY\���چ�dXhؚ��9.s/�J�7(|�:���ΤD�,'57�}�߉�(�D�d Άw��n�;j�\�����%=�ltL��+!�	
]��vz_��A:�.	���f�:�W&	&S_P�E_��7O�G���nb�+*t�b��c��j�O��]+W�
[�ӟ���X(S�)��R�D�D'*K;�$���e�J���pQ9i.��L��֍"VݧD;���l��ْa��9�s���3:V��$;�F�	]��}V+�0@=��C�`�U111)&�=1I���$>�|� �`r$��@ݜSѣ$�!v+Vl��n/��p���P�5l��Հ���J��&�?�4�		~zٲקּX�QǨ�*�d�'%a�K�~_I2Q_�x7�u��8����u��bDxv��eY�ZNey@�q011Ȟ�7��+O�X+�� ��#�0K�C^yid�:�O3�;!Q�IRe�Ø�n� ���w�8�Y��ň�;�N��$�d�s:v{��+3�ic�h�_�E��5O���g &�#5������R���BS.9���A���	+N�o{g�%�`h�l4�I��v2sv����� &ó���iT�ё��ZI"�?��$R'!LHH=*2R�ֲI���0���^��nR�%Y�Y���ΰ�$!�<�R�-w�d�R���Y_�Ðj�8^�a ���F����3Ȝ<ԟ	&�ƹ_J�
���@��`�LMI:0���o;�K��[%Q�+j��j��{�PP� �H�Fܗ����?q/S_��闖-��V�NiHMP�:I�,^�
�VK|��bZ����X ����.4ך9��}�;��%�NY���;�^�2<|͚��~�OI*�C�BW���X":�'7����`(�Wj�4��	v��R��VA2M�v>�a��2�=J��2Dn�;�e�N���&��|9�O�ݣ��/�X��h9�_�؉XJz�|ڃvG|F��pW�K{���q�.Bڜm��SĎ�0�����[/�����{|=8��լ�IJ�x:���_c��1���X�A�%;�� �[3cf�n�s�f��۸�럊;R�)�9��6�������JW�0'_�U�[�	vKs�j7�����	;rǔ5Z�뭕+���|F�zp��"�� ���g�$�Ý���JI�c@C���K=�sJ2��}w>�¿-!��T��`uZ-���up�yv�׾ƪP&dv�c�1<n4���=It�b���wP�g��w�].�6utx��f��N$1c}�ٯ�BC���l���NuLn�1�j%ܓ _��ے��q�j�$Ssqfq&��xÝbLV����ǒ�CăgLD�\�S؊�_{�ޯu��R�2��ȨȨ�����B��2���H{b��ʋ���7��3v�}�SA4��ٷo���;/��x;�2�lؙ���m������ß~����I��-�R��*5�(H	&!QL�Y(��x�]�7�����[%��s��K6o�V�h3��$H��e���w�f0���	F�gabթ����E�5���=�CB�E���8�$rRM�Y� �F�V��M�zi��+v~*�a3��I�9�jlخi�	�7�F�7vx���:��:�`X�Э���6Vhր޿����KJ��7GG1H]��R4o7')�q��]�Ve��p���s�;�+��F2�E`���A�Χ;�ld8�^Ʋ�=�n歹a���{��P�O/]�9*R���<_)T:0��M9�-���D�b����&��`��j��~�U@�W��ܱs�b���aD�s���̊�ܻj9r�ů#~���fӕ��U:�-Āq7�c#��a��3���\g$&9�>>M�[�;&Q�[��v�����c@�s����.;1,9����3$~�ʹ{��ף�T ��;�O�M78x�����=F�qOcQy����\^�]g�%�5eo����g�O���\.b�3�Ǹ޷-_��_���U�0��jU4�$���bǿ�]�nړ]��M�ii�E��E�iۛs�5�[���YɎ��-ɩ�Y��<��E�{.��z��
q��$oz��.kB�帐��p��ح�d �9�{r�>&넬V[�'�7rLBQ�#�1��R������ ��(�� vb2L.<!�]�I=�ڼ~.8����?x?��l̦Ѹu����~v������=.;��R\V!o��)���J���8�N�(%d�9���Y]�vQp̅:������9�s:���}��7�
;�,��8��e���Z6Q=�J������`O��g �A蒐�g�K��A]�^���m������;E�_Y�`�BJ=$(lm��C(����]i��[ط�lM(L�Q�<b�D!!'N,����.�3�98����UEa� ,|��o����9��/%kIj}�vSbb�ׂ}KEEQQE*WXQ��`2w������q;�����{X��/��a�������E@�N2&$l{����A�w;$�f���o�g
bBc�&c+l��)�L�YdJ��i�̽���g�<d�.9�@`�@!��#C!��*l����\L�6j��L���09Q���<_���gӲ��@ߦ��
8�9c���`wv�`{����ѱj�z����F~6CB�`��[��O&SM�Y����mN0V�3m�I'��`K �x�0�F�+v	���`��Phd5�Á��붭��}���^@��`<�>7��t|o0���є4G�J��:_�&�Z�� �{���B_���ZCM�>/o�x���E3�H��rL�����CC}�.�@���"u2���:N�����/*�tXg�.�`ys�>� ��d+�H��A֠�8�T[BE�5���dJȊ�k)�6��TA���3�������w�|V�c���3d���-Fb���/���@=��hr��Jk`��Ua�	`��Ɗ�V�u�� M��(l�"f!]�*�d�|!Z���۬��9c��g9���ѥ�1���u�:�L���r�;��B�j����Vk�I�'I_vI�*���{Ă�=f�F0��}��}مָ�x�q_c��gNK���#vLb����j�-�T��"wu�LؚG諾/X���.#yֿ4:FH4y���ykQNcv�v�a_vNNQz�#-����v�ў�\��X��dJ��.j��c�۔j�B��}YI�B���^�X�Y^�r�0LT�p��������ak#�Z-Ǔ�`I_v�ܐ�5=>�xC���d��������g�on�3�6)9.=��h�S��&ξ~��u�:���<bٱ�� \��0��5j�*�X����������1O
F�w��1_'v�{��Ap�~����4V��9D�L���V\w���,[{�B�(h�\\vff�Œ������4:�^�j����e�>�1�00v����6�%:3��ʻ�]ă�%+o2[q	Q4I&�a�%�7᚜�I�Ur�Ls�.
���z�S��6-�$�b)������؇�RGEm&�V�ww䎱#.���G�u�wJ%9�N���3�.vA�X������%�Մ�I�4TI��	&q�qIi�&ñ��ZKq����Ȁ+�~�)��t���6��iͣw'Y��Ғ ȓԌ�5�����I
�$������%H�kS� ��$�lO�ek��0�Ȋ�MB����_�*o��v����5�`
�����Ŗ�ZKIfI�b�+��J9��e"W-G������KC��G�t:��&՜(��AeUuuKˁ֦�껈7��ԧ77o5�$�Q�eL�Y	`�[dO�ر͊&���4J޲�`uLjEIq�%�b�dn�/�8p�aL5�Pj'F�X$�s�x�G��c�b�-�%S��)�Z�MmmMM��Uw�d �uOE��X�/3�d�$�_+�ӣ']sdϤ�g�(����Y��S�C��e��k�33K�2JJ��H��; o�IM6�C��m�K���w�	�_{�W�o���s�:CAB�iJ��U���h;x�pk`��-�����X�Y�Ss�]� }/�?���&�����O�8�΀]�^�g4�[3v ��ƒ���c������&ȣ�6��H���=�6�E��Hk�Ԑ�&!�2|���;Ϻi�b�h�<r��Ѯ��*�]S� ��D��w�\Z\zjZ����
�7�Y�	q�d♴�����l[�l���9�-�]�#�$�(+�<�R�5���7����lN��|�V��C�Yp�#?^�eGl��k4y���I���N�]��t��C=�u��J��A�i9��޸'k_E�>#�=�>+��㥸-[�sSYQH�ϩ(�g�u&��L��w�Ac�`[�s�3J2vd�<#���s�� 8���&���Z̛AXw\�9*��2|RR�T*��/5UU�����9�s���]u��[%SE��gu� %�ק��q�ƭfs}��7oi�b6�0���F����[g�,E^�!���1l-�P=�<���6�4�]`��.�kzx��JGZ�W�\���h�c�����B@���˨�J}�`*$|b�T%c'� V���u���������~��?|���z��y�$���l-L��V����0�={�Z�5=N2m���B}��\��h�Y�
����������.EE99����K�v�8y�U�(���0;���X��w"�/[���ea���v��D<��Or=�x�@�|�}ee��Σ�O��9�j�p��������mx�}�4XgÎ����(�"���t�$J�qs�9>����-[%þ����i����|�3P�����j��;2��3���j3��32,��L@��䮇���5�qKk}�vmf����{�/
wF��f��> ��b��ť�J���ӧO�r����vp)yKy�hHmN���������"����{ssQ�o�;D13i�A�.[2��s*�3�6#��i�cJ����Th�+W����RG��m�a���γ爖|�N�A���8s�h��a����ɝ6�`7�w�L���h����פ�D�����f�`��Z��4���x�L�6�&�[v4fe5�ւ��t��Y�:�j��U��#����x{�����=�Qjm/N��R/�*�;��9}��kh��= sG"�J��R"&.M�T����Y��a��[%P�V��`kAE��T�Da�y:�i��%;2-%�9E�.�EE�%��-�%1��^�ū�׿�2���
߃@Ⱦ8$$l3槌#�w9M��
�AU�/�S��:~�POOۈ�o�����6޹�K/�R�X��lJ�)��Ro�̅�lx���[$��9[���O�:x$�X�Vc*́�%�6�1';��6�<�ȒQ[\!bP0�;��A��Z��s��ƶUȔ�x��ˣ��L�h��nKK[�����������]�ǿ�Y�#�j���-��Vј�l�*�$Ki5�)�>!��l5�丬��t�B���4ΎOê���K�w��76e���dggזg�Y�:)�	\�>F���"K�)��ɚ��� �J�
I�Sa��
��U�����'N�qR��"�!��`�Ik��O�� 5��EY[�BANN}N�Y����gm�%Cz#dP	Ҍا˔�@b�Ԭ0�Z�r!~����l�Rb��0�;���T1�x <`_����D����0ك�|A�.� /o�j�]�U�h;Q�񑑾!��}`���'�vȖxsra|�׎�fk�$��	�	ɐ�n�7�l-�M�h�WX�3a�6���>�#ȏ�s0hD�0�f�B�^�vf6�Nc��GG���d�����[�|��A�1��6��c�;,qfFo2%�J��쥒�>�U�h;r���3�#�с��n4�1�aO@sG���!���	��5w�v,����G��`��۪��{N�=Z!b����欢�_�Ȯ-�(���@����!��!F�ZT���Va�������G ��ϖ�a���j��T�eɮ1�*�)у��b��>0r�ę�'�F�GGG��{�c�a��o;K��e�'�V6�	��=
fY�Ӟ�d��@�XO�x�eEM�����(���tzy6<���,��r�a���s���-FU�.�n'[��|���7�0d_����Un�.���e��O�I�X��:q���S��>�>����>�����N�eCKwB
�O�П���CX�C���l��'���rkKj�=j/����g�.��Cc��-i6�tz�F���6��<�`ѓ?[�RX(Χ:�2ɤ᥸�̊��\��M�Uխ흇@��;)��n ?0�w�0����]�`��$��SILK��=`�T�������eR����ؑ]Ԉ5/̐J��(�L�X��Oa2
z|p��喭i��e�&FU.�bͣ�k� �cHH0nnWk5���LL���22�Ӹ�J\'N��ltbm's�w�ot>:���؉���[�o��gd���&��Y+�98�f@�k��&�S/��f�4fg��T;�`�md�����lBю�d<n���8�N�#������}����lP��1J�ѲR"U�(
\Z��v���Mbe��^JZ��~���=]�}���_H,��U;p�w���}o*ETg��1)�<Kk����Q�����Kvy���S�^�=��kG�ϱxB���̬T��ed���*̙�C�O�Ƃ�x3$$�� SRi�"o7�X,_�X�U���p��������'O�Z�G�I�{�G���28��S�Q��� �7��g��>?	��k��%;�-�9E���j� c/dX7uOG��c���=f��Q�ݯy'F�ڵ*����=�uU"���A+�F�cb�L���H\���OڒaI7rz��������ǆ���0�q��p'��Ǽip�M��V�|�����g��b��c�ʕ]'�X2-�E�����b'uG^�������)*�O�t��'�:W�6F��Z��U����H������4(tL�ژ*1)�3���}���J6�$�Z��=m��C��F3����a� ��x��^Z��ǔ:s�j�D���w��9ҳӳ2 ?�� /�h6%�;2�u�]x��� �J����1�g���Z�NE���=���EC̎�ʮŻ��$�v�n�O*�/i�7'x[uG/����1��T�:�B9dp��T�(�g����@e�`���������-:��^��0�[���]����N�[f�8���h�	�խ'{^�c��� �x�i�Z��^�X��lbM�e+8<����md�C} �N�œ��w�0�V�c�K�ܿN��!�������F�E�������ȁ����Ȳ�!#8�yպ�c8<�GK�[��\w�-�uYHP�쑑�|Ui v̑x.uK�ěZt��>�b��N�S�8���zր�a&���,F|-��G�P����7ף���~�q:-.�Hck�~����@�:x^�s��dꜽ�����p�Ǌ��8����,
]�R� �H��N�91ÓZ d?�s��Ho;�����ؘ_�S�(��ʦ�s��a�P'dI��Y��E%�J }�IbGK�K\��K���Y����yΤѰ1j��W���۾x�P_k[�R���"ޱ�`��$Q���M.!d?�ڍ����Ї)q�����a�#y0I��ݿ6�b@�".Sf7�uKF t�1 �̭e";vήcqOS �2��hYV���1ns�����8tdJ�7G2*��{�2I�K�ǛZ�ێ�<y�Tg����G�^��n%�D���̀�㍍&��_=v!�`D���T4�Wd[��|6w�;ؙ ��9��) ;�; ���M������4���l�bR�a��d�I ؓ<&�K��B�$䵺��<}�xg;P �)y��2�a�@�y�@���F�b�YaOyN}}E�G
sE�<fZ2�1�}�M��:8����ɒV�So&�V�a5����]���kt��ɉ��g;�d<֪��6�OO����*��!;:��1Z���--��Jۜ��ڦs����3���,�b��,\,���'f/�(�L��u��_���Ɣ�Pc�XVM�=yc����/���,BŨ���`LM�1⹽���9H�CUuK{�q��N�
�vY�cc� >3�F��������ꪪٳԻ��7x�=!�|���9�>�zyvIIɎ�yl�^�=5M�t�/�� ���2�.���kB f���3,�hLH�
V O���(vO�A���;�wY�����? ����-U�����55�E@���|E.�+���Q������@�5ɂ��3�3j�{ؚ5?�Y�@�L�|Ha5:QHL�M4��ߓJ�F1CV����㝮>9SR����MՎbr��65��c�d4�5TU��t�;��&AMAvQzz}:�/q��̴�q�p��E��Y�������e^~m�ּ���cp��V�:��$Z�C{I���nu���8s���>PPf�Tc`�ݩq��-y-- ��g�*�k�N�<��9tlANv}z}c@	�[��QR����= W�fǮ����X���x'�3���}ox��(��es1<O��'b�J��h�z�����'�v�n�n��T���h ?�ZPTR�����ꦦj��h4����DF`�5�ِ�6Z����B'3@�Y".l�!�2��Qєi��kt�7q�:t=����L���x+��� �Q�Ɯ��5�קdJ^�#y�"�{��nM�)�(����*.�4_m�_v���q����z�^[�uvo���Q�Y�m�����j���2��2����0ľ9R���'y�nM��'�؛�ۻNb��u�v���>����d�jhIo�%�"�����ׂ]px��ΘU�ܜ��^��2�R��0��&�5U���9���w�a����v�(�F�
I�s9�A��,�DAjim�=�{]}Cn����̥D�CT�C�wzIIyɎ�L���Wħ���F���\�NK��T8�䴶���fB��oٔ� kK�r2,������7�O3�8V�UGo^��U,�Lۻ��΅��Z���DO܈���]�jiw�²��k���_��k�c�Ѵ�fX,�%�����Ē]�l ��%��
;��"�i�����9�vW��\Z[Լ5��6Ycg�9�^&���D�/����d�:4(hvV�c;uR�{MPm��N�<�v�oԋ�{}�X��Y;d�{,����E.�g�ݤ�l��F_vQ���&g�f��cO):�?x�zQczsVQ�ve��RwȻ��,������{̛˖-]��z\J�˿�W�Vj��0��8�#�{ծ̦CD�C�q�ɸ[Z�6ZJJr����q#v�Y�K�mO�2�W��<r"�%����������g�f7�I�)�c�:��+�q���f��i\f��'�\̃	5J���{�M��\�뀘��C��>:�c2J��z�����ꖄ�̒�z�$�|mFɎ�bx��4'��㰊����������G�����SK�|�^�]N�>��({���yn��Q�<�z=F�*\��t}𘟓U��Q�*m%����	vrIau�ȩ���c���Pyj;�wJ�4��IY���z\�A�\i��D��ͅf��;x<H��a�= Ɩ�QQ_�%�\nPZJ����ee7&0x?�]�NN`&�̶U�2�n�5U�,	B�Q�R�����jO�n�Dg��������c^�{"H�:�A6�d�Xj���k�=�qUf�(����M�Y�p�S�b�����X�AW���5�������f�
h�#66V���3:�J�s=��=��c�e�dӌJ��D��D��\WE6*%
��ޞ�������{���E���S�ޑ����ؚ�rϦ�f�t����-��Fч��b�;�N+�-ٴ����V^6�����F-�;��ny�3v��N�UEn�z�4���Oc1����*�T�f0�
b��%a�xc{)d�#�!f?����w��e��{*3�2��2-y�_A��U�]+�Gd��c�1nc�d�9��q��&<���!1��p{J���+� y5�ZeV��4'����h�ϔ�u��{�e��4k���t��S��.x�9�š���%y{���4�u��E�U.L�Nw���H�#�;�	�M�S�v:�����а�ߝ�l�()�*��j���D�YR��I6Q��6<�(�d� `Omc�:��QgG�㼞QM}zzcFV�Y)�Á�Ѱ��X�}{�a�N2�~{Js_x�Oq�cq�3J�S�񉆴��d�A���Vױ'O���Q�����G�nY�0p}���W%��Y���=���Y%Y�@�E�}�tC� "��9햒l\8-���:펁�"����p�j��k(�I6�F���s�Y�S`_��៝#3jT��A�&��;9a�����3���P�}C�G=�N͝j]�;c--թ����"o
q�D>iLOϩ�G��	v��	�1r�-,��g�`t^�t9ʟ�dZ�:������k�N2a ��uZ&J����<�bs��u�C�3U�mn�SJ[H�z�wD��ѱQ�dh03��4�q����o�N�,�eed��-(q\9��[%΄Fq'S�$8xގg�9�qEEYE��>�ZE���Y{��K0n�{��V�������r���\IN������_�؃�6G���J�R�� ����.�O���r��{x�ب���r�64��^]����$#+;C"13 ��ʌw� ��ցI��<@��tl�f����l�s��1Z�)��J�rĐ����;=�]�]��DuEX�T!$���/	�T�Z�lm7%��T�;�9���A��o����$�y�a�o�X�s`B�G��A�%���9�qxmޜ�a�j�]�fd�g!�%j��%���^���2s�"ذw��'rp:�&:r}���Le�,d��u�*F��J^�X�t�Qo�a:X;�i@��춖�>jS��j�p�v�[2�r2����gd�@]���mG2V<%������������{�:ro����F���1�@�-���b���v��S���ϽD��Dj��`UU-�Ն�ݮSd}�OY���K=34$��L�p�&HsvIqys��|�QiM}vF�`�l���y��M fx\�K�ͮ�+��� siIyEssNFV�����wy��7���DG��T!$������j!1ɖx� �Yi�n�L�Ȩ;p���������읏ϴXr*��Ar�X+'����EE۵�O,L�V�M$=����Q�Xt��^f���j�h,o6�x�W�����*p��L:+x���*�V_)��� �0�j\C=y��}  ���C�>�B�N�>H��j**.Ψ�`γ��y ����Y[��Y%�h���*J�+֘S�ϰ��uܧQԼ��(c�#�㹯�:��Ö�\QEk_ؗ��T�X~:�-�y�� �� �C����[q��!��qRu'�ŖL"k}�Q�ֱ!�ˊf�n�0���w�.Jv�=��h��P���:�lKI#Lc����W���`שT�~��r����8tq0��U*���A�����#�O�l��d2�\��Zw����=j?�.$f��e`�T^�eN%@���9�<�̙��y�/��ۅc����9>����L����+
�X[�;��2v�ӫ ;9�s��/|��/k�R��ڧĎk��؁�A{��x�N�}�z;��)��0�ALBnBq�%�BV����*�{VI��Ei�&#��Tv��"���\�Ƞ���%~KQE�{:4����`�E�y;�ۃ����>��s�W8T�<��)"���z����S.����_�v��0O���M� z7�B}�KN#��ө��~�9�O��������Q�oC��+��i�D��Ďjg�z��r��סa�1xx��^I�xF/��T��:z����I3dS*���Ro'��n�3�r$38h6H�����Y�X���r.C!�:mI���1s�Rt欌z�a�KP�^���ђ�5z��W�vF�RGn�fH��0<���Ah�k#�U�<^�y^�������Ӏ�w�c�+w�	r���㦑����0��g���
,;j�rJ�E��*��PT���*9�v$�ǝ�@�Y�>+�"\�(�gױ��hʘ{nn���ZU�f����2����dF��V�iiF���)�c��NWǨ�3l�1��T�����gJ=L��
A$���#�>����"T��2�볳9~���B�)j��9xFl	�:��]�;��]�ŠŚ�W!q_켞a�`N��������;���"Ϩ����Ҍ��ފ)*�$�K�neC�>�b�����:1�sռ�"fr22��.�}���Ɖ�l[������C�\��z���������F#��F��W;o2&��nOu,b����>�̂��xET�*�$���&�<E�Nv+�<��� ycT�򋼀�jT�ƭ�K2q�2�jqWǕ찀�@D���^��5 Cm�d�3�U�FL/)j&����3�5�-��)�#j����ǝK��]0�$D�Ր����{����_�.^��V���*Zj�\��hm�9y�L/ݣ�ޤaY�CwW����0����-nSN���K�g%��&��L �kd@xe���E���þ����,�����g��y}EQm�R���1e�JO�l��X�)�Y v����c�F���L����^��k?!��F�4*�rZ�.,��u�(��>�i��z�ST9�������%�b�h.[���c}��ͩ��./��&\1���$6����Ɗ������eէgY,q:��{�ma��;�I^V��̝Ω>����?~s�6Gk��`�)�W�����s:�F�Q��G�`�i�Q����a?<xxp��ڔ����9�VNg�=�%��윊��l+g�v�ր��	��Ā���~������-�φ����?"#���.�a�z������˛���?�����K	B	���L���F��m�n��Kw�)6j��d9�'���:���hi��,�OGΐ�=��R�Q^��c�c�L�������j�,E�=;�g6��8���5,^�9�X�����<�L�#lbez:���N�]��\�=�e�9�^s��ѿ��b�	bs$�c��@�S���{�G��i���("W��)5�n�[p�������U[��!el�j�&�����K.��d��a��`6�^�)���b2�A؍��%Ŗ��X�?͉<2��2��e����5� �<����)����� �eMZ�J�sի`�?�,1-����;�xٺ�H�7��=�m�2C>�g�F�1Y�cnR�UfT_�>���X?/��i,³E�r�2,d�V����8����l���(M�zA�2@��"��K=ò�mEcIv*�'�̈́��j� ��$S����OLF����{����O�^G���,|�����ſ:�j:�U��]�Ob��9�T�P��h̍O�b�P�T����!� .kܓ!F3����_��3F�$Ҳ$��*M�p����Q�>�)>��=f��nj|ey�0y�ePʲ��H򨿔��=vv��"i(�S=������:;-�*�~��ɓ�\�1�^���{��KL>?�|����4&C���n<�R���B�^�-��S;D!@����&�Q�>���[v�W�7♙��l,'��СeH��L��P�ye`&9X	qh�� J/������vU��M�S|�G���r_���i�^���'qs����hGx;q�����0@N�Ƣ����jG�4�x�8[\sv(�O4�I�P���Ɯ��̭^0���b$���^�S��Ƶ0��9�x�2�fJN�bs����A��qK�����z�C����
t̆=���h��|��<�菿G���fg9��3m#c����ݣ�Ì����=px�3��K��a7cUk(��������
r�n�����Vee�i��%��=;;f	O�Xkɬ́����:衂�}F��<�JU�����W��y��<�O���y!�|f�ع�<r�'b�P��}�������GF�te�Z;dK�g0Gm�nk�k�������v���[�YI���ߙ�C�~�l�7�Z�+j���ir��3|�N_,�YE�8<deZc�J9�&�gf�LzNI��F��Rp�����]o;SRR��/�}1%%OvsxM��,0$a�����sf윎s��T9���?����Е0�j��tjǪG;�pkۑ����)����\�>���><�ɜ:k�� M6��&om̐��p/'^Qd�c6O�2��hڊ��fgz�^�XQ�c)*�h�*�m?��&��r�÷.:a������=O�z��Kix��yy��3U���sy��wu|�Qo_��/�R���UQx+���UMq�iu{��gN��uw���:xt?6���y��`�H��������,`p&�1U��,p�1���F�����JD��d���Xo0�kۂ���/i̪�.����U}Qf�YC�e�:o�SR �G�@��?���) r�~����7߮S�c�SR`��D9��䶾���peyxM�O9	_��kr���_�I�G�ɲU�dK����S�Q1~<6�7�؏�:�r��������}.���,�����t�����l_�V<���>�O�Ɋ�9Y���a��}�4��f���lxh%%ȚrjK����ܱ�T���q��~�Z_�����Y�✸��g�Z�ݹ�.*
��7��j2vR���k�gp�b}����=�>Ŏ�Ah�PI.�n%�vȌvw�z���9;�9�s�tboo��t�&%���T�_�6���9>琵�<�"�ڢT��d2L��S��
KQ}V�%Ò	)RNI�����b'�P]
��t��Ṉ�=��t�C�\א�?��K���m;#����u�RF��)��s,��+Ŏ�z����K?��7_B��Q*�+H+0� �'��������%���j�m���9C��wv���m�;<<08<-�����]��(^��'��xH�-
7dgě�iz�"nT2q�%����l�1�(Φ��3愝p'&�ч�c S���y���ߋp:7�w���w���7O�{���?��O�����u2vr���f�ш&S�+���(c���^z)8(,_�Ҕ���nߎk��[Z{I ���9�u���u���1l nw?x�ȡ�Gz]�Q���T��Y���m��g�k,/W���۽�3,x�]��A�i8��D	�D�h���qcv�>�ۧ�s�M�~�����1�������{��߿0>���ׯ^����������`B��;b��UUJK-(HKK��ؑ�W�
$IS|��o����pĮ5	|�d2�&c�&�; ��~�h穃m� ��]��c���t�����ɜ%����������Y�ob�]�����4ؕC�y��i�Y���bɨ�i�A�z;Ω�kW/]z���3��SRnNDL\���{�㗮\�4�3��~�xO�#u�4��A@kװ�
�'�?�#}|��o��/�k"5���d|Uդ"$�~��5�v�#mOu8Q̱�m##�G����<c�}z���B�
BI`��=E�`-X|�<��v�Q0���n�b�NDg��ȩ�.�)в��}Ŕ�DN�׮�������;L��|������L\�|aܙ?��r�_���1�aȡ�ʨ������b[�y�)�R��\L'c?}�����Q�@�b�<��;r`=����G{��Z���;��VO��Jn���`0w76�d�E��ۦ�n�[�p��Ĥ��gg6�bxP�<�2�)�׮^�z������cq���w�s&޽|	xG���������w�اS;���ޥJ�S�'c���~����/�G�4G�=,&�Qi�"�z-6k`!���i;t�s�Xϱޞ�##����Б�Ǐ=z��1W7]қ.�A���*yLFo����۱&\��3���Ѧ\��a��zN/�ygKy�����k>�<z��+�\�p"�!�G����իW?F�vg���O�^�����}���&�)^���!0�Y�D�:�g��y��D���r�ςV��G/��,[�U�!�[��W�p*�G��Wǀ��Α��3@�����遠����#]}�'rZ��a�;��WskEQ9�/v�D�[rE����1�(�r��6N�P��+7&�]?���޻|��k� v4��3��W�^����[uX��0�`gx^���p�΁?�`��/|�{?	o�,c�����4��&�6I��B�su�\������u��{{<��^�G����f���^=#v	q�T��Q�]o�L�/v"x�HDC��|O�8�I�ktvn��TCi�R�M��@�~>�}�b�ҕw=��?w���Sa�Q�"���&���4��A���=�@E�O~�lz��*��ռ��^c��V���9������(b�Ԩ���c#9�r���w9p��($�~%�� ���ψ��	�qOIv��̛�ԎA>�fP���0+�Y�kt�6��.c�z�F��҇�+��.S�W.�����~f�|̗����;p�%�Mk.�Y&=�-+�ru`y�
��'��%��G���/��'����R\�/{LUIR�F� �D2Gz�@�mX@���#802��>0<860�ڇ��NcY�Ӷc)F�|�`5a<i���L~��bv��m��U�G�1L?�t~�>
<⣫��/\�~	XC$���f�]��|�!N������b`�
~cg5س�7�yM�����,	&�uI�6[�iK��q˖}E;2�L�l2U���{7�6䦇n��>��q��:
������m;~��{00[
P�,�i�*�JFI4H~�`&�����<?����tJR|�؝���M��ML|������/�w��K"���7a"�s{��}*��\���>nKsFq���Fh)�W=���O��V��n���Jv腴��=��~ݏڍ��p��PG����> A��:�������~vv�6��6�.o��q���'D��(�=:wg��W�u��;Zp648�!9��a\����g��|�>L��|�����.6wJ�i��x�&��c)O�@l#���P�=�����&�v�W�KⰌ��S�h4	��w=M��ݣ��������Vױ㐮�����9r�Xo��{tpxxZ�Ӱ}V�(╜�d3��˼��� v�;�g0��a����Է��%���G�}��އ�}4q�\~Jp?��{������?O�N/c=��a�:mAFF��&Q쫖/}�!���c��\�jgq5�eg&�R�eG�)�9�%��~�>���E�������>�.w�nw�Z��[���3��e�;���\o�� Y%�����{7`9��!`���w��<�6�,���0�m�q8SR��Md ����ss�S`�k��I'0ƌ���vU���xi�{���쎴ڒ��$G�}kq��J��������h%gj���h����ݭ��qlzo?;x��2�SaG�cc��� y����qp�]����I�F.G�A�y)L
��<��ф+אT�P�^�����
�V�`iLƊ�F��b��oz��ړ�J
�JQ`�g� ��x�r7v���1(���7Hޡ�On7�?�;D.12u"xr���Σy�o;f��<M ��oLW��v<�sa�\ցO#67w����)���q�+Ț+�����졲�)� /�Jcc�>�B}f��T5����2w�y|&�C��j��c�d5�q����d%�������T��I]��&v=����������<2���\:��\���M�x�gغ�1�"�q0��}��Q{0b�i��`�S��^XW�#3�XU���G亯r.����7��~��O�����F��I�� HD쒨���w`���W�l2��t����g����{@���?�����7�cE�w�����H((..ά�ax:U{x�j��bw�Y��;v����`�����N�����C5��׌���g�>�5VWO{I�L�m;��(��e츂v���Y��ݝ�v�G�uD���~BX�����P���t�d-�Q�F1�Փ��o���=����-{���d���Kh�cc>��*zp�lj���l%j���fg
��p.�҇��.������u�2�6�+���y�v�~��\N �a��>K�A�; �V=��	v\���iiU����ۇ�ce�=VC���`�7ټ@��`�w���`2ۨ�%�#66O"���L%s,��Fj��Ρ��e�(��s��a2�?�#~�����{�j��ݮ��3��wQ�G����'o��bW��yV'���������~R��?:0�=4pv�3FG����F�ãÃ�C�q�;�6�=|xxԇ=�]��;���<�I���s���@L��Qӏ|R]
�����PQ�"`�P�sl�^9�2��>���54���N�8���g�q���a(���Ù�V�� ������cض�L�*okq�Y�d�����@dL��Ç��vHR��e�>mo:<t�����>���>;I��Ó��+VJ�#Ȕy���w���@"v=��ΒԐ���/�L^|��p���dN���'�)�H#H2���Lzm����\n���^���.{����|�C �������Ѩ,s(q�k �c�>�1<�w`���sdd�p����9��� <
r��0v�>�[�L&j�"���N�1R" O2��;�N _1111ܝ�Έ��Ⱥ�F���!Ź1[f��R��#�'��%��;�;��<[�rL���x^Χcuto�G�?~3(�W�1+�q���K�vE��b��nW�ѣG��FF��:�s���j�<v���#���>������] ��>W��#������ui�j7I&�� ⅊&��{��8��W�o���^~;�����&6�w^8��e��3��G�ރ�������Ͻ�ߌȯ��h��}�s5��xQ�3��Q��~�e4��|s�gJ	����=�EŖ4pz�`��:�����}�;��x��k�����PωC]##�<t���h��С���Z��\]�r���d ��ҹ�#'Ox̻A"��)�
L`n�~�*��y��_�����/�_8���˗�xnb�һׯ^�o��x�:|��n�ElR�<�t��z;���:D�<c,*�lܷ��b��Y�n�E=ϔ:�R�M��X2�3�˷x��j'��ɱl������Bꡮή���:����TOO��@ϑ����>W�уGz��L�`/��~��II�ȍ���R�1���<p/]�z��`�ɥ�^�~i�����.�x��{�\�r��G}���K�>��~�3b�������gg�����;�-9iH�ױ��?��샽P	������=�r�is�M����u��i<r���C����ރ�n��1|}�T������[1zv��KoO�`3� 򱱼������X���*]w"���W�Mܸ|�Z���+�o��/_��������O�~2��y��CP��%l$HI���O��a�1�IϩO�b�% ��������*�=*J�g����oG�]�1r��k�ءS�;H�h'�?��{�(5�S�}ǻ��Cm��1W�CgzG�q�a��݂������&�DFxl�,���{��XRdt�����_�h����7"�/]�z$���E���#���<�e_��� j�1H�b�0/�1@�4]�#�)��~�cĎ���4�v\��˹���;�*8v��q�^wG{�3m������;�{���v�F�69�3#]'������~��2vyN���1�!Bnd�0z�|�δN����ץ\�0د�� ����߅_'b��r���: �o8�/|H�S�;&�T����9xZ-m�]�m�~���:�����W��]�N�S��!������\��.l�C��hm�<��!��؇�G�Μ9����:��>xG�E<������:���EE叏����'�P��.���ꕫr�]j�/\&&���K�}�ʯ�/W*��V��a�Gƾ" {��U���Ԯ��P���~��ў��3��``"�#�t����{�xOϱN�dd���ԙ�'����i����;x;�B�������ŗ\���S�'&O�č+W?��:���ĵ�W>�".\�~����~�����TZph�Z��j��}�c��O#v�FԽSmd7�B��`?��������=�sj��,L���_X����8}�>ꃹ�`�ņ�1!���`�����_:��а����<(����ODD8/]���ᗯ�{��'W�^��ة���Sq�o��;�
[�Ț��&��%����.�h�^Mz �w�F��1�\������?x�Վ��zO�9�s��ox������؉��zێ�8zx w_c���Ig[揽�j-���5����LF�g���f��������4u���`(W�گ_�v�껗6_�����?B었�{�����ϐ쌎�`�b�埅�(j���R��OJL�q+�ɶ<'��@��=]�C�]����>�.W'�����$	"���S=�!�9y� q��JU�v�CN+q��9�Иq�y�G��#j��� S�{����!~����oL�����`-�ǉ��G�	;�q,�c�=�L���z���L�n	�c�g4&�UV"v���m�;���������dr�6���C��`v9�$n�S���|��]~A��M���Y��;=�T_װF]J�\xs^���̿u��ȇ0��`=��<"v�گώݔ�f4�D+�}������0ȑ2~j����%��]c��u�Ads����=�C�M�͑�;���T���`�qu���~�b��N�.�1��<��E���(�.���E�|]��w?<�l8��yV��]�
�a�4��j��2�BrAnJ20:V�N.h^��G?~	���)9وeU<ʇ̪��F�WVWc7�ɮ��C��Ly��!l�=�;�կ�#�����㮁���;2��Q�����V\F���9J���"�x��{]�͛�����:>�����#P;`���=b���/D��� �y��3��U�d�~;�~�;
z��l�9�����{�,xx͛�S��@�W�S�@P�9��&���n��}��u�9ER�����vWVtº��F��<0r��qrP�azf��A�`u�PU)ν�?�b��v��Bb
�����WQ�����k�3pt�R!v�(��ĥ��l�>��>qr(g�]Q����X���X���Z�2vߚ7�ՁH�^V��.W�TY�Vx#���'1p�>�	���!R
;s��Xױ����ڰ46���1�v�O���Y@��v�T�[�;�����w�ةǤ���<�ʵ�n|t)����� k�~	ˎ�ͫ � I��=�sHb!�G�z��c�X�7�����V��#v�;��D\]�N�[�3� ;��h_w�����<t���$�j`�{��A�C�~�ࡃ��v��&�;Q{K�0/�`2(v�K��w�=7��.e�^엯^�wi���������Ό�.I���o`�tYç���a��������l���޻���0<���*��g��ޓ�U�}l`�����w��������2ǡSxK���:v�H[d�mG񡴍�9+�1�yb��]�z^�*���&9Hn�3)���o8?���+Wpo̹	�k��x�8��y�c|s�G����k�7�G�{����H�~V�84دA��߻�o.&�`g��^Ew�@��ݣ�}}í�}�7}}�Q�n�B�!\�;<6�doo[/d���a�d��yc���:�J�Ǝb�C����G\�t�¥`
��>�p:oE�GL\�01�1#��"ƣ �t�O���<���ӎ&���_��u�́{=�؃�6F�� ��i���cCز18z�@��`.`���3Zq�}��P�mo8{vpp�E&ܳ2��A�����N:�~�`e���N��k����nmw����6�㪩�y�aW>�j��4��E�p9�XJ�:?***�aW=��>v=������ytip��b��ㅝ�I(���=8�:��va�{h�o��������qxltxx�\P0t������!��vj2�2|�ܱ����n/c����߿���+r�b��~kí�n����ٰ��[�v5��������x�� �N���Rx���|騙v�VUG�p����ȗ�d�VF�u��U�t&S�O�;	�"}��
,ߦ7@�Æ�n0��N��p"U�V�ag��x�U)-�<h�T�����}�b�]�c�7?P� �pf����E�Ȧ`����O!���u�n��IS�:9PFE�EY��Cߐ6Y؟]�Җ	BҔ� �֮�'�w�t�Q��N����o�;H�Ӿ_z�5j|H�c�ʧl�=놄�S��M �q}�ٯ?��3r������
�|ٻ��Ex��".���ŋ�z���f��hj�wO��y\���ʟ�`ϴ�ϳ~x͏�Ɩ<P��d��ZUZ݊wG���py����Q�zN���>�}H��;<��o�w�J�֖g�.����e|��/~���B�:���R����q����I~ �����yx����6/��Ǟ���2��y_YM�f�65v�����9l���Fa����w�Bp34�׫v��"�v���gϚ�9c���s�ؖ>������7(2��6�>���'�o�o��0�y�{��59#vž�H�~����F��j�F�����NO�"���#.�e��ǃg�������A�y��ym�jN�%r�8v5���׿��׷���ߥ4��%Ö�Oܼ�ط�̫�n�R\f�b�����@{�]ܴ�"�����⮦�:�;	;]���_VǪ��
��o����~�$xq6����&Q�t7GUu��$�{����.���c}�ۇ�����thЫv�i�0'o���H���Q������v��8;�,��r��3���]AԎ����N�N�ב�M-��S*���ԋ֎�V!v��$���K�����F���d���˩G{]��}2t�r-��(�f�J����N��õԽ���P�JKg�N���-�������ǮoصK:z��	��-����]�<Љ��??�Nfٍ7��}��Ι ���)"��5�J�B�}�s�ޢ'C���%���GF�e��%�Y���;}�t��=J��Ue<�	��& ;���Ç�j<�n��vQ@�ča�������0�}�._K����̥@�G\��������7lڴi#�N�?��ѥ�HWs�c/J<����N�j�c }n�X������2�0�$�٘��j�<�Vw�Aso�C����&�Gq��'�T�P{���B��Bz7f�nC���.Ȳ�dF�`?;ޱJ�=��l��1����=FV;�E�.��o�$؝޽z�	g���%��f{��`2��Z9��{'ʂ���ž9J����lOM3K�@�IX�Ē;vt�(rL~����= �|+��:9?��`��-�!%0�G���>���·��:�A��������#�#�Z;��e���w ���W?�������@� �Ӫ�d��K"����7	����6���$�Qi�{u{!{���	oB�.����D�s�-��>[�Ύj�ݿ��/>��s��=��=FQ���-%h��~���j���<1��k�~��'MN�v4�Pe6�j5����}��xd6�����V11\[���$�I���N�SO��v�tzgĴ&3i�F6C�����ٰ�;�>#3*��;���k/�>AJ�^�[�$Տ�E��c���'_~����)��'��ec;���g=7�,X��7C������V�`�$g'��]x�����n��#�1�>F��)��Tj��l��jr3Ŵ�����ޮ��-��w��M��co�+x�j�I�N�ԛ�����|ą�����%�P�S6'seM:z�Ux�j�wi�����Qb�<3�Ҫ~W`?��+v��þ���j�1�A�Ui���r�V���A��s�2n��:L�>���X�M���;�b3�e���ҕ/?�x���ع&n#־�9��n>����\��Q�2�������{bH�8�;ih�D�>L
h3�Q�g�*��q���Χ���G��d������o1F	e�1$1
��'Y�N}�S�7 �k_��;s�e���zY��]zdF����5?��@�Z��M�=�4�.ut��ǰF&�1���6��ٽ�_�4�����M�
���A\�kG���g-UnѨK�$���l����	e��v��Oo8q�4عP�;��G}/�\��'�	^�.2R��D�Tح��������S##}c���tN�z��iG6y�pf*�(�|���$K��a�=]�\c'M��w�l�-=�����/��7����c.�J}����ey�V��;��|���Z0�o��#,�-���U�d���^ZU�\T�G���v?�ϊݣv|�@���*
ʲ�����G~�{�~\ǫ���~�g���������Z���Q�e\�;x]*�x��o�b�s���
��V���a���2'��1e�Ri$3/������w�+�V�|j�ݏ�?�ˏǜ���$��0OK҄���1���S��i����O���^5�D},�G�ku�(�|��>����������ᜪ��S`��i��>r���\��d���X`�8�IN�{�~v��A�W)xZ������?�UV�\MF.��}��}��$�2���� �o|�)�1�r(G�_6�2-�����}���v��/�E��q�x� �U�����<}��@��ȤJ�%?���l2���`uu<���=����א�~Fv��U��U�W�c��^���`O�vE���%{��q����O�r���A�DΙ�v4���ýAx��6τ�ɯ�/v+d��--؁z�k��T}��%Y�j�U�T���5T󸇇��Ҋ�(x�uP�dA/��䜱��1��n�ZO���؏��3���8x̧�^r�9�����}�^�Nf���-�Ǿ���~�#\O��I�elD��.�SiË�;\�zN�<�َ�逬v9���ۇ��vy����d�7��E�*����m�F��
>?��x���S��f��~��d|B�@������x?�d�G��2j,Ȭ\��v�����wC�<�w�jY��YM��;�B^�Bz�Nw���r���\n�#�1_��Y����5x�oKuU����`�Ng�X�0șֻ<�z�=M!�^��@���d<ޮ���$u�	ڱ؎jϝ;$ӌN-� h�h�O��CHp˔V���xCAr��W��[;����k����do�T!}U>��'ѧ���v�L��;�פR��Ɖx������y>��/�X�^M�͚x���1������w�ң�6�KK��>>N
W/9�p�~j�ds�0����۰3��@k'���-}�i\a���$^2��lO5�c�A|'����N�&�i�G��>�i��;YeR� ���aϦIeK�[������v��3����nrZr�T����2�ڽS��F�$��%�1uux:���8l5iF����hz��OA��?��ݥϐ��:�Δ���P`4H�&C�%[K;ޭw������}�7nT^���u��g��&��{�`u���w��˛A�>׈�陙�F�𢡊���g������N���O��;1R
pv�$c���A.d���@��y�w��5@k#�1ZC���s�Sa�n��N�ːUo����~&��E�@�l�]�`��"vR~$�'�]�v�:���E���#�9��E�{�\���U�/�\�0�.6 ����q���̑���ǳ�֎��k^ziiHв�*�Fc�E�7|��?�|eu�������-��J���Y�䒘�ڇ�6���n������M�������Ϯh�uXr�55t_�nݜ;��-��,s�ˢ��	��qg������.=F���֯[��k-��}��_�ђ�����[�x>�4	;r� {K���Ҧ�GZO���j�,�'{�'_=|u�ė�W�*��~�E��f���b���ޛ{o�.E�ɐ��e�`>N���c����;$w���e苝D�+V|�{&c��w�C����H�'�b v�H�x�[{ۉ�'�t�C��r�>O���Czվ��������N�ܫ�����y3aw(�))NB}���N���o�Y���}:�$I��A8�B�Boϛ�:�n���+���ES`_�̩�K����Vi���j��'U�`R=�L��{��[{�>m	rF�z�g��5�:�5�5�������eyv�}�O���a(��h*�+�w�d��{%>~�/]j��� �+7�x�>�ڱ)�G�\����_\0���	��,���*̝IJ=P�I�QF6�>���Ak��$����L�PF����-�>{�����\y�E ��y��2�모lJ��|J�ap���i3�J��?�I�q��`�|�����/F�y��R��ؕ��5W�1+��Y�����{|ُ�,	��pW��R~�,EX�[{�b�:���x��'[���ˤ��;2'[��|SH�yX���.���=�0�~�~G������}��7x[�f��G�����/��)P�LJ�WnD4����~��� ��Xxy���=�.{i)�=|"?*Zǐ�]Id;�w��N�>�4wӦ0Zq��}n��`�W���M�A7���<I�> �x�:b��;�ӧ���z�TiЈ���]&��2����j|?�
v~�H��1`17����*<9�I��u�u����/�y�ŅSb_�0�� wHT�� w���J�`L�kj*q"��fΜ�:�«ǩ�(y�s�x��A���Vdg8���o�?�ݏ�=�����C���)�[����&-�n�N�t�	�'�,���(yˏ0�b��˫7�	vR~�˵z;{����W�~��gL���[M\f��H��Q��-[ s����O3]=gN�9�=}�}�����(����.O������f�-wZ����b�ͥ��2r^�B/s �����D��8y�VcH��@�{q����$���ٯ\�"X�r̻/r\�����{�-���NIBH�2K�����K��D:�^
�#]�jj�`�
�C�q����R����a�=f(����)���ᡳ����Qse��*��>�:<���B�̚fR;�(f׭����V۝��|���k��:}��g�b�C�u�l�x��M����-]�.���j��|����.��n?FRՑ�Q�@���l.��E�Oatxz�b'���L�������Y0�ݿ��{Y,�G�N!B���o�<�����n����֮p��:��S����D��wN�ؿ�ri<?��s�Ɇr=F�s0�&:v۪W�C��ӇN�}ያC���F�4ح{2OL���=xd��?գ��a���5���>4�ک�鮨Q��u��w����<)/����B����c��a�b޸m`J�ߤ��S��N��<o�������:��b��b��,�4�sժWI��i��G�P틉�u�d�l&�a4T�D�I؅�k�����@�G;]c���c2�:���gM�hql��PLwF���ݿ��琣b������S���B�w)�(����J��7�~��������E|o�i�<������k���o��/ u}��ỚG�J���9��]��R{��o<;�؉ˬ	Y�4�GD���Mؐe((L3�;aH$��$����1,D�(&#����n�8r�n�a�9GfNj�����o?��n���L�%��8̚{)Zm�0Փ@oǍ�����������/ೆ��"H��5r�a.�k��R���F����׿�b�t*q�gWä�ر�W��VsABB�YJ�}�{+����!QrӮ�1o ���Mfx��i���[ �i��5����ݿ����|00����=�NI�c��>���OV�u���jG����FV76�^��L�ݘZ�j�Y=`W� ����E�c_p�#k����Eb�)��p{������+�6��{ ���qTn!��.o��_m����?gT}�e�����|���e�X�t���j�r����wm��$�5��������q'����Tl��@���2�����<�ң{�e���b��7A�t��g㒪�巧�M�ye�ɐM$v�`�{�UOg�w�U����Y�.���1�o�u ���o?�=04�u��Q��o*���w���>�}q�L�`�8y����7E�O|B��$U�Q�o��;�-��
�޶jU���ן]4=t"�ܟ!whYS)6n �Jk vR}�nu���=5�F�c�4W�������.����~?����w���v���v���?ڰ7�d��i-斢v�c6a�43v�r�%o\%	�+�aG���@�z�x������r)�!՜VcÐ�jK���o��o���UU�݇�e����Q�2Y�S���b���X;ʽ���| �F��ü��iT~s\�E�  d?IDATj買�j��췦Î�#����vԺrbu v̗X�\:�ry�˫_��3b_pϓ߅�i�3a�j�N[J��&cG�1	խ��Po���=�v���f�9�}�{���W��X?̨_�~7�;���cS�!�wz�/��0��7��X��j�b�v�S��0,��N���k���m�W��X3�"j@0s��!�}q��HuLG���,xXM����r�5�-�-�m='Ϝ85�k��ݽݿ>U�)��Sj}l��a����8����L�&�Dƾa���8�*�I�6���,j'U�M�n��OƝu�!=^�1�9�(P��L�u�1ʡ3p�瑧�B@&U���^)J"oc��{23R!kii��μӽ#}l(��f�o���\��;�����ݿ�fT��Ô*c��9K����Rk��X�/��T'����~��#�ƹ����1���K��ix��Z>Ky�	U��}O���ZVi��Qp�ƭ%��f��Zh���w�ę�]�c���crmfxlԷ9'������0j��8�z�JĎy�D��L���o��U;Q����=����p�XN+��Xr�31ϕ��#�!zT���.�;6̄,�
��(�:�n�9�D�||��b��������u/18�~ػ�c@V�'��jR�
;���W�`��l������ީ���}�-n��[�Ș��}�8̧c1&%E�jMq������s�)��m�c���M7�y�VP�Q*MYUi�++M�����zKN�wWWc+j�����'{���t8@jWc���:���ϡ6�F&�M�z�NVk���ۛC(j�0��oFx�\��oӣ<|�{s�)��"Ĉ�4��d2ec�{,E�N���Ife��Z�b0UZ�M�s;]S����ݒ,�'��$)����qO�e��u�*SUUu�n[KG���O�< |�a��@����͎��7U��A�h7$K��-�� ž��d��ME���.���6�o�!;���Ť4q�Dm�5[���U�hc�c�_ �S�N�s���a��I� �G�"�Iʄr�D�6�紕�+U��1�A�LU$��Md͐ChP����Ge�˻'瀽���7A���i�n����>��}&�+�r˛"�S�>���kjH?��^�β�4`�j��ѕ���}��u�Ͽ���9a_x��T�e�4%-�W�u���L��Ί31�������R��������'N��(��D��u��46;���?��ގ&9���X��}���������v��4Wu'V�b6���<=�Fy�O�Ƽ��(��kĮ�ë�uQ�/]�s��,��].���Hș�y��P�`�j�2��C���M4��mխ��Ev�ww�ݞ����/̦e�I���j�'�J��c�n�,�3�/!~��v��
�~3_��F �MX�o;���1���z�n��䝾i���ȸ/s�>C��ry)*�J�m����3��<�&���׃˨TB��3�9;2�tA�l�\`����@/.4��J$����e��5��$�#v�>�o��ݻ�7&K�䁒j���i�S�D�^o�7΂?n�bop�'�Ӏ֯A��%;��66b�TH��<�J�Jٹ��_ú�\&�o�����j��I��p���4����$c��J<���ڎI�ɮ�v�I��x��V���pr�Xw�,u��%�_k�&���{���"<f�]!>'�$}E�7l�0>~��_^�60=����}��>oWѰ	E%i�\FGZ����+��{�b�����e!�zLU5�
Kc*�ЛL�Upxk3���ʖv�"O�i;Ї�z�YS�ڇW
P;��OA���~�G<�O)Oi2>��6��Dl�qK��y�ž��y�����0�+�^p�1z��)v>W��
��6Ƹ�$c����3�%<�[s;Y�~=tY0Ye��o�1#s��!k���)s
^ �$�<�7v�����B�l�,���!7=����?*������`2�������:t��x��v��#�/��"6��}}ľiR�2����;↙�7"���i���J�k�!y\LYZNI���E�m�Mb�?w��NU��ɐ��Ie��O�D� T�Cu|�N61&
��d��4r'L�ȎU7�I��o<=��nqv�+�i�2�ʥ����_�����0h�@�`�uk���4������3c�8��6l8��޻/�I=���#��x�#b��26�O�Hž�_��}hќ�c�C��!��0�j���(`���rD��PY������G;���C:��	y��Q��]~��ݯ(]!��	�~�����HtI����~��M�y�X�]6�!N���#�Ms�NOa�o���2�~|!�.�6s�ەK x��(9��h;{����n1D��[B{7�GF1ZM��O�N��*!1�z��k���S�ǈؑ����v��!E��!�b�����[&�h�;���w��}�,�[S�qS1���7����h}��&0lGj�����=���1����3������>��C���y������iY�T�[��ƀ;H�bUuu�ȡ�3�O��ã����tہ2��}��1Y�C��tt{_�&F쾻c�$KP�����{ ���z��'iq�wD�~�dGr����CnE������_�Νu���b0>������<���M�떿��s�,���}쩥X ^���F�k���N�c7D���Lo;p��b']K�}7:�1?U���b2݄s���_����|��P_���e�Q��%��9���~+@�3b'Ա��q'9A<ej�d�)��v"���y�]YfZ�) ����+��C��[���8y�x/6��̱w�H�wO�?w�c���j���88r��=��Q����`gY�h&֓��q��f�T�.z��f��r2�q��x���w����{-���G�R�"7�ؗ��6w�Y��w���_	��u��Sb�[>�Y��7��u���P�r ��	�����
J'��Iٍ�G)��ݿ��s�ڻ�口�j��M�"1��Q�T~����kױ�q"��\j�B�i�����%�i��:����[츚M��<��j4�Lv�*C&U�j� ~ {����*�U��zzN��떹+'[ ��
�ܣ�S�x�vyA�z��1J��RQ���~�bQ��i�!e�t�Φ�7D�_�J�b�u��<�/W��+���sH�w0�QEm[�n�߱�����B��aV��(�*c����.��c�w���By�t��ҠG_	�)�k���&CfO� /��j���dKk��c�4��m���e�؁�ƈ�@�ˏ�͔�L���;n�F�@I�s�	��=��7����7�}$(xɒg�Ƴ}4�;�H��h����^���F�)T�n�zS�N���H}�|D쿑�����M<«v�P&b6aD�;�zk�j���󘣮�8w�n�p6 nl��#��d�`�%����X�3�n��#9��v���'�`&l}�J��$�m�UU���/v+���Z2U������q�����P��T���e�S�����@��H����[���T��o��/⻈�dez����+���#"n\���������T/{�����؍5&�!&���*U���������~�#��X�	Z�6*���L�`�k2�%Q�De�oΩII�RiK+V	ΜD�[>��ɧ���&V����7�����>p��-y �2�z�`�6�m�7.��i��צ���I! '�q�8��^��%��|܏+��&�>CwY3���C� �aYV���u���ϡIcz���DP0�"����2&�LJ�)0�@�|���1k5��{'��z�xg{w_G��zT���� �O1�v�	S7��ݐ,v�|�CM�N�Gr]�����e|c�&N��;#n����x~S��=Wt���!p:.�f�	��!�|��u�f�g��ܟ
��=w�E���\��,�u
�I���]�j9�y�����wR'P���q?�ܧ�����g	�|��P��P; ߶����_�4�M�ȈKW>%��A�y��s������h���ֽ����n�b�Xx��AX�]d�њ��`��`2����JB�Wwp�y����wNU�>����dL00j��7�wW�ʫ�[�j�HՎ&3_�+?��6Ab��׀� �qd3�$�۪�hX-��Q̊Go�bȸ�ᧂ{0C��њR���e��tTVUW��$<�����>��'�Y�c�n�W~�����縎���ңv"�m$~$זȝ]�6��d��N�q^t�ߠP���	T>�);���8LVN˱�,����z��-��̽�|78��"I|$q�t��X)T7��=���ޑv�1�}-{�7��q#^�>`+k�{5 G��OĎ���ݷ�c���yuv�yܐ��~�&�l�%�s��^���8�V�0X��t>+y�`_��O�%���m��ju�\�J}�WS޳�Q$��x��iO�W"�̽o@��r?�wt{���Ψ��o�Z���I���N���&���4G����$7�
�������V���q�&K`@}�L������
�c�Rt�:��J�����n�����~
��#]#�C�"��,���=@��Ed>�sT��O��Y�dN���ۥ>o��rK�x�KȒn����W����;��ƎUP$�s��	_��F	l2���^�t��కQ��*'*���$A�W��Х�*r~5�qp��nwɗ�*�=F�@����]�ߍ|?�;���d��5J���2��p���z������o��x~���xo�Z���駟@nZ���v�s}��q�T��������k�-_���7�~:-������JA��##�:�\�ѻ$�D��e�0�+�;�O<q�����j��{`T�NW�����;|� ��m��?�����8���������6^�I���t���Ѐ�鼘R�0>qm��O&�Ν|n�G/�D�z�J�O��i?�yx���u��~�ݰ�{Q�1k
'wjx=����I����l�3�&~_�z�X�Ϝ�lw��:�;.w�r`���^�˓���x���݀�H"��Q;́�6m�6e��̩��+w<�g/8�0y��	g>��NOn��<)��ȝ�{�ξ��޺� ��y�#�6=������r���e�*E�dlVA���ɍ�D�粁Rwk{�A,��mo��]��(�O�>_t�j�����G0���.�F<n�[7/"�%t�5����q���qD�3%������m�H�2'�#_��5v�uu�N�b��P����P���Qd�J�cx�vI`i&^������%��3mG�;�q���2�nxvc	��u:�S�Go��Kl���c��Vx��U�Q7)���xo���p��y��y[C����^����H�M��� >�ߟ�ϓ�s�"kJ�8�s;��37�_���Ͽvw,�p_�����d�++�F��LOMƚ���dR��K��2�a�M�t?Fs�X灎a��F� ����N���D� ��>�@������8T�.�op��ڴweD�R��'��q�u\6����;��Ԕ\�Γ��:r6ΰ��&��1P_���+^q���3������b#Wit�P�u����n�b�j���ӕ�w"I4S]��ڇ;�O�8��NO�%jw�
2oA��cH_�w�+
|����׿T�78�:��^=JNׄ�O��߰i)�*���)���В�T�ĉ��`f�����z�G��\>V ����^Xca����p%�D���C���{okmcZ��mM�BWl�T����\���iHـ'S��a[*dN=���ۻ=z�|
boQ���]�z7b��]1��-g�M-8�������UW���z�!roM�"�i��S�e����A�GD\�v�.V�G�1z����<>�=m&��0�XS�w�p�\*0��h���M���puh)F���f�U�!79��%)Q���J.-�"ۤ*ڄ��&5��='O�tu"x�H��vw#_4��~E_|���<���bZ$���$+�����ݢ�������������rk�ܧKσ����Q�o�?�ĸ�K��QT��f;]~!�x�#c�^S��5Z�J�g�~;oooz�����5�3��C��V25#$$;x���&�Z}��o�����>��!�<��jo���jmU�}�Lzv��������j���g'4��ݪ�����������R��
�u45v�GJ���s�Y�0���?���/�)��:	 e�˟Ô��݆�U�;qi#�����q���f�g�EFE�5�i�/����=��L�R/UIh�y��==d��݅�b��--���>���䨿F����
k����d�m�I-JS����V���ܛ�+��)Mf�r�o�̆���`.�����&�lgR��\��.�2Le�#F�RE�\��6���!�\��sEB��{���H�|�^%�$��[�-I��tWwt�<u�4p?��:�>:8@������'�Q�����v�������|_Ӂ��_���MM�����Kٕ�Ƿ�>z��6R����=,�nڸy�����W>�4�D���v��WĎi*��XF�7Y�t�����r���W�YJ�Ga�w�-����RE� qb3�����p;��s�Pϩޑv�pwk�B�bX������樻�t��t65���&�W�ꖦ�􆺆����5�`o�%_�����~���q\9�|�y?�N�0uX^�u�k�;�iF��<LSIGu$	b�V<�û�'�'5`�V�`Z��ְZV���kܴ�U{��[J&Q�L����hN�siW��[0zA����pF���v�Êi�nښ�����)-'^�PW�����?��'���ie��x�N�$C��
��y�f�w�Ong��̨xь����,vg@���w�'}�1�y��eX{���u,6�xB��jC����+<�dJʓZ:���L��'���hom���0n�P;<�Vl:��g���w��DSS��Ƣ�&wK^acj]CC
����_�S��@�v��o��[��tbԈ��O.��ӻ��q��^��v=$��H���5�ߍj�4��}n�2��g�Y�ʩ��5Z�F_IVY�6/�J)w���:X
n�=~��I�\�9r�@��ޕOZ���j�Mg�V�dF��-M�%�y-�`��)uu����?��D�B�����8����:x��6����K�/��(��9"uދA�N���,	Ӥ������XzmM��%tm�U�J�j1Q�$A����+���5���y�P*�hW�P|k?�d�g[q
�������������Eg�~��_5�@�[s��>-�����&y��dS�{��7b)~�N'V`��H���9���d ;6�����v�ZC�r� �;������}ѳ�=�z_BΛQ��ʪ�$<^�q�5f�l) _j#)UY|{{_ס��Ϝ>y��E)�hW���� =�̨�zS����&<��������T��z;�sYɸ��z�ۅA�j���q��Opķ_~r	�/���Uw�m�t�/6� U���<���
 �U�+捯�:n�x��5�h�J�&���
W;l��P�f�ԕ��0"�7ADS�v7u��9y�oCţ��tx��z�{5>'9j?�3��r ���Z�nii��hL��P��VG�U���*Y��}��g
�w��L�(��qlqd��zsc�aP�!� ��b�k< \��ڹm�ZܢԿ:���{)��΄;����j
���^�����1@URށ��#=�O�9q�x�Z���t�z-�7=r�/���1ԦjwuSK|��nWC���`���?���{�>�'?Ҁ��1R���+�.`���er'a��;71Vgޞ�{�ɱ�jr?�u�.���ʩ�ߋ�>O�3�A��]�j�d�	�&��"�#uH�$�NV�t{�n;�s�s�L���ʝzJ+9��3�v�ݖ���B�6���W�bRv���q�ڀ�?����7�!��9�@bF�H?����%g�����X=#LBN�N��'�P���<8�:ZA�[�;����G�g�g��]��hy�h,��@�B��D�Dp@�WK��ɪ2A`�R���t��=g�!��ݴ8FF}K��ϰ�q7�>�kI��quUSSAcӰ+e���!&1���vz�TyFG���NfW'^�g�����O?�v����Аߠ�\a*�+zs�ɜ���rh0*u�N���][ś�=�=
�*�����괜	��M��$���$���TUﮮn2���e`:�h��1b���w�o�WC���5��q�_��qk�j��Rv����?�k���ە﹎]��qܣv�^
a�Eg�s�Ƶ�����0O�y����|�tj��3��5&Y-b�� �	[������T�����k�]�x(�����N*I% ����D��ک����yeeǃՌ�?M�Q"����ؑ��_�3�2�"��ƌڒ���_YҚ��S��h���oc%̩�����J�>>N݅Z:��x~T
��I�b�ϰ�$�z�����l&���w�ĭ2+��.l����ױ#iV�UZ]���MK��f�R)`f��۳#�)C���%��׀��|;�����o��di7����Φ�MKN�,�W9f<��.�����d�kp:����;�m�$bw��4z����?�v)������H��ܢgrqC���91���m3yy:�V�QGGt�������L�����ax�_��22
������Yj�A�.��!{9멌��w��:t��ɟjs8@�(Z���̨�޿�m�/B���UK�YwK
.*��GGE��5 c��Q�Vs�<N���O�G�"+�zz~J���>��^��e&���cEN��u�Ѣ�G��t����1M���C�����K�<�W!wF�V�b�Q�]�ٷd�=w(�Q|{۩�(yȢN���P�0v�3�n��2�����xGJJk
��)Q���3zcْ���[HQ����I�ӫW>�!cJ
�N�]1,L�[�����b����^vVYB$�z��_/u��R��WO�u�|�Ϊ�x��� %O�Φ�na��;����4�i��"@�ٜ�"��nv��5١'/���η�cI�%/%'I��c������Fwc�o:t�	^Ў:�z�d��r�2Q:���y�5���O4�&C��1��m=u�G8�4�;���C�τ,]�9
^'� t�
<��!�&L2[z�����_��z��'zͷ���^���n÷(���-/����Adiĭ��&F��#7��\������On\�p�q�)�?��C���wyl|I،�o5�5�|�v�S�\J��&p{ҋ_�l���^�
K�|s$&�}R� XMb)�HN0b�l)��|��mخ�4!x�^���A՟��a�m�=nkojwu�y^�,S���п��:/�=����3���}��2����r`"��]F��P�yzN��*8���b���KJ_<�'JG��֭%M�/���Sa�t��?
��A�-_��c�zQ�؍	Ɏ@��F�Ô�G/;e@�`�h6��C'Im���3GN}����n?@G�R-#�SKKK?��� \�f'Y)�'�ŉ�K�ʉ�?�z��sh.0����P�v���f���/f̵����sx;�%�}���~-Y�ܟ��^ q$YoڌI\� ���ћ6�fi_m��qǱ��� 0����v��)�Б�v�:~�-G�����<�N,\���'&@�(�+W�
�?�#���+�Q�x�@ڻ^�k*���;�Ʋ�#O:{�%���'֑Ť?���@�.�%�P�� ^��d򶧚���`�[�5����p��G��ήcG���9��o����9~���Q@́��|'��=q�*���?��Be�)X˥��|\¨����\�(�W|*�cx���e9J�L�D8�	&_�h�Z��y�:���?�P�S�������%�8�(L���7l7���݊]�|V�Qcwp� ��8k��y|^��JفvWoש#G>���#=$�!�s�����O�:v���^��/��q�І��*�nNя����R����2a�?Ƌ��;�=%�Z;��=�;.($N�թT�h�O��'�N�?�E(i�|&��̗�&���	&��b7�8<{d'a�;H��~| ���K�~�����ԑ�'it)��4�=y�P����\�F�p��y�ƥ���Kuu��X{����ƙ�+�ر��R��F�B_ߌ�#@_�'�.��k��,�y���j�fQ�L4��J
v����'�㡸S`��w�G�z�PE����Nk_oױS��P��T�ç'�F޽���N�r��o q���Hx�9��+�)��q݈gJ
}M&S�(�Z̑��v������ů9\�<.z臯�YBN����Ԍ��'�K�i�]�D!!#�J����;� ����E�h�r�>�������sں`v=
N��s�>y�ı��W}qB$�ǀƉw���zn�;�b�����[ �9�6F�=H�I���𕏾��V�U����Р��� x��g�q��O��\Ccc'J�O����y�~L�e����|F�q��i6������u�رS�#]����҅�h�$H�C3gR�w�����ә9<VWPR��D/u�^�;50Z_���X��_O�w6� �}~Y���g/]A��B4�r0��%mٱ=�A}�����1��(�o���Vr�8�N.e��^�8�@��]Hܞ��'���c�9�No����i��;��?Q���X;�0@$��:������p�k��������SA���}HF��V�TY�r�v���Qae�d�$��#x�dZu�1���/�w�(��8���G�XSS�
�JEґ����W0r����x4��͕�O#���bgD]MI����i@hł�DS�gݺ�嫟{�τ:r�y��χ���h ����hbtn �j�XaI����?�y����U?��^8��)z y$��<��g���j`rC0��|e�r��<o������񞙖��ͅ�.WN9��m_`둛����V�jܾc�=�=�|�+�?�7�,^�����1��� ��ĕ�s��9�<�epb�v� �c���Ho����ȳÏz��_��Z���s�Xw��y.7���&R�a�t�
����e��_�s�NR�G���}q�����)11V�U铤R�\T!0�0=v��'��<��Ͽ�5`υ��H>�j^A��Ǆ�pW.D��2�=���l��?�����s��mk��W�����]��X������g�y�o^	���1-&��ccKKM{2�X�h��n�r(bW���g`2x��jed��h3�������}��@��	�0�j�p��(���;�	[��6���X�}�/��Y�ʊu���?l����j����f&�g�+�(��`s�~��W�ӏ��?��/�c�!��O�$��V2�%�U;����D��]��>5#�L� ������ȑ:
��-V�g,X��#O�D��Jx���?l��DC�ӕA~����5�`��s�4��^����~�먟�^�j/k�Wջְ%'sGqF}�]�z�1�}��;���K�1���+7����!'"��Ӥ)��{y�G�߼����ݿ'�AΊW����CS�L}��S$f�<�g�
&cW��/+�qa�eGfIfIqQ��ȅy����f��\p+����,F#��?���B�����?G���$`_����_�������֪mx��F��2�<��?R%��;�KgT�QI������x� &_`)�I3'o)/�"��%0��	���"�INx��c��j!��1��\�v��|�b�����״�!؁��,~u�������=*J��@�id&ўÑ�f���Γo{�v;9���1�2>�9�2�������&�ݛ�����V�w�%{��'�t;�K�N
a�1�����Z�`�����߿����'Tľ�ľ�#�������?W��DGk5��2v�pw��6�v;K��+;��@S���!�yj.r�^V��d�wץe6Wb�DԞ�G}v�����+� �L��8�:��hYr�������?�tJ�����?�����c��}���r������/�\�j3ݩ��&��<��0<�U?Z�gh��9Įx:���ʶZ�r�t�A L},�>�ڱ����9��L,�_,���uo��?��m�Q����؃��oP��c��հ������V-_����;a� (�������i�v�*��˓�ˮ.��+�bIא�/F��c�+�}:��<f�?Eҋf���T*���j����x+R������<���b����g��!�|�{���?����a��?��oǨb�ZG����q������	���#_L����b/S��vr*��̭�����4K���g?�����^�5I ��5���ڶ��ۿ�31�����'�<�B���3�2���"����?���W^}u�/����L��ߏ5KX�ϵ�v>-�[[�#��k��N�N�\�����LKIq���:9�7	;������̏:�/F��T�R��`ԉ�����������:����b��W�m�i]y���$��I�{��U!{��w?L�U�/r��BH����%�%Y�i[=Y	@������3/���$)sw��o����3dqbs�ַ���������.S��2��4m���	����,Y�A�g��K�й�O������e���k2����������m }�����:�-����H�?�k��op%�;�9?l�����>^�F�sS�����x�>�c�?@�e�v��UVm���6�v�fytc����� \졓/�.���p��cz`����/��ܾ���/ɓ�ۥ�c:-���<���/��/�>���"ۑ�׏�Ĵ�Hu�:���v�U�]�B��7����i9����,ti�]q�b���cA�C]�B��te�R�Q��\[���/�,l�%Q�S����kd����~limka�nOY�a4��Q��5p,`vf>0��gjͦfRU���a��q���ˆ'&$�w3�����6�D �4,���~c"u��$���d}�����z�N!�%�J+�v�H���N~e��Pjy}��k�+"���j,��g�k���__-CwJ������G��-�~Naw���x��3��,c�������vW�#��+�伻��ď������1�>/��m�za��+��+~��/8t��ߍ��&�!���8�e�`��A 	t�A�Sln|��~c�y_A}�G �lB�Z'c�Y�V=+ 3mK����	�!|ǭ�>�1k�y��"¾�{E����P��	2L���Nپ���x|!���b�����.%�ޝm,�w��[��_�^���u�x�8��fE�h�H��ޟ��`�K�+�n7_5�LcjV�����X�������[���l��xl���n���E���ט/�_]Sy7�E��U]k��vB�sK��[kbYH�/��|rc��Q��;`+8CK`fn��^b'���H>:��)�z'%�{`�}Qj������N�,��8�D����Xp.�Lƒ[�y�&���㯩�V0��vd�x-���?��{�]���/vz��E������%؃��/���r|+Z��������y���5s#�z|��e_B�IP�.�_a�"��j��n`���j��`�Y�\���7O�g�$��z�χ�͗�ǘ~{�I�F�_��P��%��m�:?=�w�D G��v_���v7��tR�8�P�_�Ç�vNK�n9\/�s�jWa��ۇ�u�w��ɨ X�j�пzҎ�������g}�.�3~�`0@�l ��`0��za���t���.�ܻws���(/����� *%�Kj>���~6��%��<�?>>�����P/]APm�oدٯ�&&D;CH�{�&˘Z`������;̅����.��
�N'��B�g��쒱Jf��f:�/<{�Q�qH���3����g'�E�����\Ӟ�$����l�a`�"v���z� �n1�6�49ˣ?ʾ����ڼov��[>?Ĭ����@=#!�7.�;q
�j��7P��c����"/ ����NC�s����b�n�8Ie�8�����3�Wu��Ln<)@fxAg���dL�[���]�=0���&b[k�[_��t���/��%����_m)R	���Σ/�&b;s����q�=nTcRu�[�}����F/�'�eDe\k4YAfxV=��g���< <@�^�mn-�����B�� �_ �� ���Q̇6ׂ�3��,������5�8w�7�`w��_ߎ�Hv�U� ��4�,f�]5ii/��� Q���B�eQ�_�4����������w@���^`��dr:�)�yx��-��\(t|�k���/��8�"��Է�Kv$;FL��"�q��d1�<�`�s���:��_`a�R0��>C��/�.��#ޢL�HZ/��5رj����!?�=H�	`_ �O]���&�Z��#�)�|]��W��rE���0�H����8vt3�,zw�B����ւ�������/�������A���S=0����Nd �P�=�Nʷ6d_�M��6�P�����2��}
�(2Hw*��ĻC���>_�-�e���uB�������`��LGv�l�_f{൰��!R�vw+�*��mBT��ߝ����q��
�n��)��q2}
��w�#�d\�H̄hg@�Y�j��Y��z��$����������W���5�h�����>�1�gQWz���G����f20. � ����+Н�ǵS`]���E�%�������vd;Uw9)�;z�U�
BUg}����� %{`e+ء���`�u\�Ի�'��/ZJ� �D ����`�,}P���o�8NW�v�dg�W�)����K�~�ۧ�E؝.ަǠ��qk�߿x`�?�Z�xǙ�׳�/ҝ���%�/��@H�S�܃��P��L�!��M�o�3Н�s����A�A����ò�������^��pb������ll��h0hO:�${���w*�bf�%�g�9$�H���Q�~��	�}�e�rY���B�Z�<ٝ�#d��S<�������z�Z�	�$�(�A.��2æM��� � �<���\2�=Z3;3�)��wF\p���l,��2� ��
7�u�%;�z�>��l��#]�>�!;I�qb�jġwV��s�>���!P�5��H�ގ�e�i�zѩ��� Յ���g�=��#��_X�}sөZ�����F��vp�ɮ�/�"�N����/I���EZ�,�)Zſ ������t0iL�� ���I�Ǳ��U�{M�+5P����Z� ���P�f�Ou��_Wt��02��v�^��ܒ��9b
~���J�L�弦t)vpG%�.����}�����j��뾀/��V�g��R�} ��T��%yvb�Q^��^�'����䝷92NfX��1P��	/
�b�&��&�5�����?�������e���K� Na��]*$3��:��YÅ����Y��r3w<�I0�u'�������
�PA���A�1�����dn��j{5z{ɹ�8{�����O�x-�~�L��zaG벀)I�@,�}mk!p#Ӯy)٫�ĸ�|N'�ҿ{��!�qr��N��r9�N� �M��ɳ�z�ZԤY�o���|`��}FD��/:�)���{�L��>R��������vz�Cv��M�����I�d����А(�7ۭV��Q�)�<~z��a�-&�:c�� ���|�#�?@a�����;d!��fAD�1>���oacef}���a�hcD��]��˙�F��l�k9���ާ*C`��vk��p�5���@��H�H�n�Լ�v$�����.���I�&���/��Df�hT�.x+�j,�n��ndkSS�s�N�e�t��?���p�f0N��ק����d`Tn��\*EË�H$ф�Z%�ӡ�њL�lŲ_��������@����kL�;i��YO����%����Y�+��tfc�]��J�r��lBk�2@�����vd�|Tg�:��&B,F"�p4�l�Ԡ4<15.�wK#S+ߘn�V�fz�N����t���ɨK��K���n���Ƿuwy+[_X���������:���Z�^�;Iml���m�ݬc ����t�a�5��j�E#��������͝�b��hW8�;�Xu1<�{��i��_��^��D�&a�맗��}��<Uw�r�Q��|��/�=@�ӭ��?pm��̱(�G��Ԁz��w�I���9/�k�&�����3;�R$zk��p��WwJ�B���A���11K���V)f�����d��.���%��Z�8��ґn��8.\�u�����'x�>��B����(sk����H�OYl7k�œ�����p�� �����r�����H�o�o��h鼦�x�8N�;p�Zi�׻:�(�	�Htffn��W^���.f����@����Cԧ}Ӵ%�����}���g���g/7�"yͤ�R�]�F����{��oo�;���#����o}
���+c�Y�F��>8�M����y���Ё]P��MM�ƻz�u&J&C���?n������}�N�J3Jӗq��4PZd;W@�?�=y���\���o����������ꔪ��.�ho�Ñ}��o�ܼ�F���k��+�W�y����B���|�m<Ӷ��^j��.ir��n躴V�ŬY]]���L� �G� �����{������2�:��f`/��	\=��8�������}���>}�tY�i�צ�7���C�дn�>܏&�m��{��>]���;?��϶��ޣ�6�탳S�ݬ�$�v+�WՙL{lC%�Mm��c���V([�|vГ):�.�������+��z�rx���������'�_|������?��o�y��ӧ��cq�:fcv�0;7��FJXsxp�Tk�s����_a���D�� >���C��x>�~�CaW�	���&S�b����㨙@۶���}���������מ ��s�$���3u�/P�i��<	/.|O����Çx����?w��o�ԏI����ƸlJs;�X�١:~r����r�f��3�&�ܾ�Bp�l?�wx�Ӭ��;f�18	�[�&���Aa��.�{���b	=���|�	�=Ca�(��'O_l�b-By�M/���G���vT=C�.���ʑ[��Pm�r��-���{��} yOTv����[GvW"�N��`6��!���p����x|%��l��C��Ӈ�o�*#s�y��3�t ���|��ɳ��>|�b��J,����?��{$�������a���m��%�+6�{�]N�v�oaaOi�� q��ۇw�m-���R�4�����	m���|���L>}�����9H���<��A�����)v��?\�x�����ʓ 8�ߢ�y����{`��p|�9��U�S�]׬�E$�S�S��D#e�������qz=e��NI�I�Ʉر:y�B�м`l�jU���3�%���7�Qƀ�1�z�ŋ��i|��8ay��!�����P�㻡�o�7���>==}��i�'O����G�\�ft1"u��#�;�H��ǰ��^�y������쌓L81
2�b��	���i���X��V�IYX^XX__�ZX[��ڂ>v����5�7���t�$��D�J��xr�+%������K���w�kǫ��^\@�	�;恹��vy� 
�(3"��@(ҷ�_A؛��[m���R؝N���#ٝ�V�I2mo�)�wrj
���o~s�CD���������C�����ut|�L���
j�<t
˱/�����7�D��"�Y�lm��x�9�=��K��Y!Z��/�	�;j{ⴇ�T�B7v=|7��H���=��I�����y�M ���������<��ק��哽�T��ƃ����6ԏ��1�^]̀������t�zt���WV��@��5�pfQomܾ-х^�Cmo���_����Wboډ��G�?m����1�I��k��<3��]!d���@ڼ� �؋��- |j�SX���D�i��&_S �t-�:��z=�iu:�+���H$\˂�쬠��M~�`�
g���G��x��B�ۇG�H��ϰ�G���a��Ы��G��^+���V�ҰB�O6�� i�6���c�_��;��TRe�U�QV*S�z�x���j�Lz�m	<�ګ�GJ�p8Zn����S�tGݤF��Qpq:0�᯶:��{�7�H�������qT�1���dp�(Ѯ���qK�N�� ��V 2
�Qfphإ���7��x��U� �l�F�ozƭ���Q��sC��	l�W%g��"d4*dG�\��9^^η�f�e���h7��9��:L&���x�=��0¾w� Q*W�}�/���<���t� �i�=+��89ưvK�e���ƍ�p�H���� ??�&[H2���/ܽ�x������&���j��h��[���)��;�i2�|�4o���Q����qh5c��qR�׏;-�W�~䰚̂�3�ˋ�3"�8 �������~�]�3��D÷�5��ͳD�����.c��>�V��J^�����:�3,S*��L L��V���X=�?�m�"x��:ZPv�A�2�0���qF;�O�m��]�q-8IM�
FS�]���-+����lo��"�-&�N���r4|<9< �C�zpk'��\���a�l�`o�"w�g�X���Q���jf�dGN�F���dI� p09<A��N7�>��*��ʆQ4�I�p�}�7���,�q^ʛ���:�ł2f1�˥�77������հ��z�W���`�ZL���b�����v���w�&���T�+����ص�~����k����<)�߼�"���]���r̫s��&�3��!��a�6�5pJ�AOf��gy��XJ�M�6�bW��_���9Z��FA�-����������=R� ���>�F��1
'�pZp2PG���
^��m��8 N�<8;J$Jm3N��+�3ާ׮�vh�H��8=:M@�mT�h�Z{ݞo@�:�>y�K�dh�,�qtqr��� ��8�/����( Q�����A�q	����j�Y���@-��9��U���6�12q$|*��[�gi4Z�,����9������&�
:^\���j�H�p�sz�HDKGG�rP�W؉�|<0zM�o�8n�4q~�l�r9�N� �߂�ު9� u����dl��mTg�8���y�_A��9����7���� ��6��^Od�X�F^��4F7fjd��f�a���D��4	�&;N��d��0fէ�z�|�9���ެ��h�P*%JMG���������O��3�qh�5,�\Q��3̄�
�X-�J��h�Lc����ao��(ׁ�&ӧ��*�!�g�R�+9��Cԉ�w�@�LPO�J^�����M�v>[);�D�ť<{��n��-;J;���5-��M��k$A�q���`��xj6����>r�*�f^���zs9�ZN�A@J���o���[͜�2vm��v�li�7����0��
���[p4A�i��Z�Ly�:\�M���j2c���!"$P�F��R�V�M,���L:����Vi��bj�Y�nxl�
��,��ͦ��n��9�����!Y?��/?�ߒ�n#i��7�3�!�`6��z�"3*�}H���зU��}
��q~��S�b�����:f9�L�f>��6��"۩�d�VS�R)������N���`dʙU����
f���a��{�YPH�s<Pz,Z�R�#�>f�� ;.}�N���	�����/ʃ6�W��V݀Ld; �hۖ��ޮYLf����qM%QG�� �a9��V \W(���p�ި�Ou'��\?�o�h����,�T����Ѭٍ:'~���m4M�1�0d4R&���H��{'�d�-�?E�q�$��
X��M�Ĩ�r�շ,�r���+��_&f�4،Z�b�9(�:�;��5���'4u�Qu]���%�>��`t:l'����"�n@)
��0'�5������ZLz���Ŝ�pXA���Lv�ޟ��o����?#k�	�@dr�(��.��&�i��ㇰv0L��mS;�N��"�K.��z �^��#����;WB��h6��Q��l�` ѝ�j�k=���@���C��f�k��[�*C��hX��?�� 겫�;a�{��9��`�V⁣m��y�Q��3r���縜ծV� up1.�j0�V�{�S���8��xN�h������T*�` ��v�l�{��t�uf���w�Np��t	Qo=��
��N��%vH��@�>f��?�Lڢm�r�+3��-���(���J��1�v��	#c��`����lY@�͐jdĄ7�����v���x%�w �f9���q��`m5����jI�K�I#�5� �>]J+�N�N ��Yd(�W���~B�������U��s�9�q�l�-7�M5-�ɤ�N\Y͞�[M�l��E'cs�ɀ���a�x�jYM�d�lg��b���k5�t�ARn45�d���v�1C[�6Z�q�	q�D�K�h{߳]����I�"��=$�2�i�ZE�RN�v�#�ɚK��E ����Ll�bXM����L�b�ۇ5� 쵶��Ơ�.�C��ڋ�: G��'��q��Q�U�O�0u`�3�nBl��\g�8e�(2������W�#�.>�]q�h�[f�q��ݨ��K H4��ÛM ;�w�"�C��3�˹r�ba��:Q��R�b�Q�B�{	H���0�2�[���7��#&�('�"�0X��fp������Ô�����������hq!���R[L$�錗�f�u�k9�f�	\Nf`��-�C��r	v�v9��z�f�����M!4�Հ��{��+4�SD/c���X��m��2ƿv�~T�>f{/�!�6�r˘O�F�"���Cb��83���:Dl"9 ��n���#�l���b�煴f�?��� �� ����13j���N>�1ٵ^3<ILs1F��:K jӣ��Tn~$l��5�v��ղ!M�k'�-	iW+F���z��Vu�KΝN�
��\.�7��J��c5�u�R'8'$��Or1׳�߃�r��T`�%���A�dH��A2�@�x�ѭ�zlٍ�G���'�d}�9]N^�+�]\��\�����*���ӆD�j�U�4tN��	��C	^�}�/���d��3�I��'r��9ḙ��1;=O� ���dc�l��`�/mpB$��= �!�(���!ꕏ�qv�#�����
ժ��$�n|8�v�˥�u^�l]�&��؞ča��Ni{$R�
�	o��@��r�����.���"s��D��P�;q�ԉ�q�b��8j�Tug�Os�P$ΠB�)a�c&Nf����>C":M���^D���|���'��pd+_c�b���vُ��͓z�.���*��ள�70n��Ad9�P�U ��;���ͦ�>P!�i|�[�ҋ�7w����,c���CBl	l\��v�\'lw��L�\�,a��W������kaP��RU�8����E��rst:��ɮ ����
'�aU��0���T4e�@�	��M8I��>���DI'+HV7#���6�����T����p�$U����X�Lwg<iL �#q�V4^�:�-jW=,�DJ.�U�P�iY���Ҍ�Ө�ǒ�]A��NVU�ZP��6̠a$R#��7�Qk�P3��w9m$݆8(�b�.=N��Q�$�,EͱU��!������480�k�qD�n�"�z\/ST{=U�R��i �� h�j�G%0Tz���Z�֨9�F7Ó�Z�?Ϥ�&+��""�� �/�E8�T$_�e�w�R	-
��I516o�ެ��xF6[nZu�����X�ޅ}��w�����ҹJ�,St�9�&�4|�l6����ʆ�In���K�1�L�֪UU9k��JW����*��姨Oz��t&ϧ�V�,���8�������8�;4��r�V�TrY(�r�lת8�=�K���l`�]����F*l�bp���Z1��TmN����o��f��L�U٠�D���k��&�N�z�ڬS���6��?W=Z]���i��PW'5�r~ey!��g�^H:���zl3 %^�"��3��Z��݈g�i�(��b��1R��۩����A����$2�`W ��b��}G^��j��Ф��z�$���3�lE�l1����V��{3��բڃ9�6~R�kf@�J*�Y�d�^MYm��������nl%�O�Nz0Y�$p�� '��|<� _�43ٍT
>U6E�&���%ܻN�Oa�Ba~	w�R��r�[_UN��p4*nsA7��������F��M��@L\�[�Ҕ�G�V�d�W3j�$8��\)��v���p&�]!�)�WS+D»��ӣH<��Y�e2�f*4�I���T#�K��ޞL-E"���l<|P��hi�����_�vИt%�����Lde�O�� rr�p���l:_.j0��GS>=+����Z<�5��<*�>^+Ď�N�T�]��%�&3ͽ�x���<Q8�W���W��M�L,���w���h��W�8J���2����N)���[d�yN���s�M�=�/�.�l��V"���i�<_<;Ϧ'v�G�ΆCK�R�]��*^�ɷ�N6U:-E��T�ݬ�f�l,<#�?ɮ��@9�މDV�l��|%�����(�v���TznhOfu&�N�K�h"z�:?�s�Ψ������b���l�S��ZK&F.k���.�)�?y�K�I�s�H$M�wON�N�E� �T.�YI�"�r%�ʕ�Ō�,{�Q>�-GO��p>�h�pE��Ug*{'�Bd1�G�@jv�1P���x�T�D��JV�W�eB��X,�( �S�h���{:���b�B8�l��e�E���~iLƭ�!��sc2�4�2��aXu&[Y�$J�0~�hEc��5yi��T��(�Sة�2^��Tu�Q:.��\-�sI`O��+�p���6���v���ŕ��H�.G��D�T�trce�$)���,�sjĮ���L|%�� �w���������0���}�{&l��m�_1�rH���v���$R��Tބ�?�@�]�
 2`���qW��ˍ���p�4����^���A3Hg㡕0Pwo�b�HDԧ����N�,��2�^��G��R�di1]�zZZ�q.`���l� �S�{������ᗍ��j������;ru�U��Ef��T%������^hi/������V�P(�
��<���
t�E����04�t��ھw���>�~$� ��+'�dv7���TY��^�	o�|�;I�EOR{�EB=���8�Q�h�P8?�9:�Me�F�R�qzәh�b�{{'K���e��.��y����7�B�/K��a�U�#x��-��uv�<��3�$NRU�S����n�d��d&=������b9_޹���V-���LR�<�b�qg����ݕ�|",8�z��v�p��(|�Mm�y�VqH��7�<$����/ ��d��p����ݍ���G���;j����1 ��qy	x���A��N��[����(���L�<�O�Xu��y�����՜��;y����d*p��!���%�`�=*M�V۹u�<���J��Ȁ����k�ӳ[ �WU��x�K�;g7�����c��ƻx�������I��9;�[��R�IMV}%\y����ܴ���XF�1_��� �Qk3��ӳ�����՜���V�a�b�U�4�l:��70�� ݳ�|��U�POO�Y��<�\����O%C��w�qk^�&]�T�瓩�X�[0�8�k�lQpr%���U�.��g��r��ͽPlwc��r��D�]��?��o�Ǎ�?y%`��qT&�	e0��׬�sG�Ȫ�"8�x>�M��^���y\��V�4bE��d�0�*T����\�0*Vk.g�7w�~������#���}�2��e�MN��M7�M�PJ��d>�:g^!�v�a�2��{��1�2o���#���+d8�%�9���Y,f�O0�dV�V��nT����q��Us8 	gWFb�gFD5�N��U�<�@fh
\7�}�#��Gjĭ���V�5�|AȔ��%��"�\�4j����$�����!���c����OFF^e�U�VyV�q�Zɲ�YW�d2�8�e[�$��'d}���%y<E�	�l�&rA��Jǥ� ���n�M ,������/�,��d��VCw �j©-WU���x�~�p������tU�L�|��~ݍP����?���Q�e��CC��0*��/ޥRO�#X�<�n��q-1���Y�K�󂖡��8�zy�*Q�Z"�Xi�5JI�P��l�]$��Tmdn��_�(�*Y.��ǏA���>8���_�ݿd������g##CC����~r����fP6�Xˆ�ޏe28��Q��`02Y5@�U�@�:�3�~�0@6��p�uE����>�|i�*�pQ� /�x?���W.�����$�O����ݷ���Bt���>�l�P8��|��g�	���O�򡡡��O?�����O?��׆_�?���C� �8A�& ��
�OȽ����g��xdp�VT�#�?��c��?2�R`+3�c}`e��n� �LA��2}��{�~��[��5�	�?y筿��>"e��k����Q�сQa�B� <�n�j��1��G6��T
J�w !e�>O�/×#�@0�w���6 �1��7���C@y�������+/2�������{����!@��7�;�w�z��i�9|���ﾇ�ny����=���^z�{:G��K/���RyW��P�B����;o�A�w���x/P�S��ƛo��S(?O?��X��g���wb���=pK��gx��n!�wJ�e;�y�W
}
-���Dx��_���\�ɏ ��)�bt�r�G����7�򕗞A��y�+��9*]_�����d���1��   %tEXtdate:create 2024-04-25T05:12:37+00:00�L0B   %tEXtdate:modify 2024-04-25T05:12:37+00:00���   (tEXtdate:timestamp 2024-04-25T05:12:55+00:00����    IEND�B`�PK
     ���Z�����  ��  /   images/2abdabbf-059f-44b6-b68f-d45f0cb3c7dc.png�PNG

   IHDR  v  �   �;ߎ  �PLTEGpLT�?,Y��󼽽)9HX���/0J�D��r4��M�����*������bcc=Q='g�'Zt��-+/E<a�i����VT���#AB�fP��2q�����G889It==���C|%d�Q��<�����e^*������#VS�---T��)Ii���:) x��Ef!"Ey0k��(I���1J-�ۇq�%SUW..2���Rpsst ���V�Փ�����Av�0��&A ]�966��55#~�#8d�c�zud�M,cw���/D)�����oC68Z��6R1�����FFG���Bo�]����9X��!$��j��[�&q���ǫ�\{���b� 86	"""5f3h!fo�R\o��~r��#&"������=;���t�4M1O<5A��>Tl���9w�
00*K ���aNFb�����_2$n�බ�T�{��&r��TIA��C��Wz�#1 64(Wx=pSg��qo���";]�����O~
r�Y"@[*C&;Z111���	ebfhkp��#"IG99>?@���%a�9��h�c�����ꛫ��R�1o���q��v������*q}�������M���m�\\]@MMN��&*(`y+uqj��������! )3&zz{������%<!H0!mmo5Q0�ŷ~>�B   �tRNS ������������L��Μ���������������ą#���������z������������������������������������������������I������]�^����*���������������������������������g�����������������������7��������������������������������
����������������������������2�    	pHYs  �  ��+   %tEXtdate:create 2024-04-25T05:12:37+00:00�L0B   %tEXtdate:modify 2024-04-25T05:12:37+00:00���   (tEXtdate:timestamp 2024-04-25T05:12:55+00:00����  �SIDATx�콏s��6�F��P'&�vH ��3N:�ȳ�N��k@�/^1v�y�g\R%�pH<x�;~?��'U�M��;hPɐ
O'�k�Y�kQu�� �׌�V�Z�b���x����ծ$c�6�c�eY��K׹����>��0~?���hjj¿M���?x$�=�������-6�l4���osPď� �+~��n�qB�`��W��G����x�����W�P���민���/������'�X�O��>���?���C�!��~�5�#8�ho�������Ga�>����������
���>R��_}4���/>|����}�w�{ｫt �G��~���O6oރ{~	����O�v|��A��o:�/<zK����.�_���;�^��zu�ի�<����	����W�t ��w��p	��C�R����AQ�!��;���/oMOo�`���o�3���[x�R��v���߫�����ىp)�Op���<1��
@�������MhJ�!B�옘~k���:�Fss�N��޵��w|s~�ٵ��w�le��
��A�������DG'`�$����1(��/@V��ߚ>:�����5�{�vtt�y' ��رc�8Zq�~�?8vl׮�� /Q'����8�&����t�L"��g�}����H�=Ӕ��W;�F�w\<���9jM��Tkj(J��O!���{��_9D�
��̓/E�����r3<9 �����e�@��h�Y�[{� 9������	�#���(��"�8��l�x��ڷ��-���� ��mh(Ԋ����wp��7���K��fZ45����9L�}�;�(
#y+�����2�8�α�0��0l�-��(�!��/��qҥ�������Z�S��'s����飝����@r8
F�54D�k����6�����j���SS�=S�8��m@D�H�H��[���s��}\�N伎��o���'߁t�*˞�Np*�>�q<5���l)�p."	�*��Q<D�ŠכN ��Ӌ#�n�(0���@���C�(�m!.�8���.d}/B�z�6�0���?�@]P\z��5ا�����U���X�B ��Xd� x���g��N��t:�C��<<Г ��*Ώ"����7O%8��Q���="��o��ΈΌ�������k��Р��� m@�À�e��k�B`�Bʻ�AJ"I� d�$d��ԏ��	AzR�h�}��3�Ԣ�=���������A��C*�h�����!�*�������yExU`�.$�PHH" �S����@R�i��J !�nI���R��J�Jq
�(�D:նο}��>B�?�, ��Jy�]��*��=��6C@	�r�x��9Ni>�T4��W��XB� +=�`���^o�-��wI�����x}�ʍ�����E �+>4t����;�aU�͓��"�w�O3m���[�� �B� �Ā�����JxfB��6|�S��y×�mv�|���
T�*<�VT��}p��2��"��m~џs������t��t`{�_��7�A�E�7o���w��W�4�3_\$�C��G���T!���^��-p �t�..T	*/ �Y��r�S��/�%^{�ༀ����AU(d�>�������?�Fƿrg�!�Q�����_|��4ӗ���ڝ(�`]B!���S�
h��<�? ��J�L5�}�s'�;�E�#���q
�e��G�偿}��K�1;�w���R���\>��߂��]�
o>`�W������ӏ�@�!:���t��s!q�_|Y^�a�(p�'��at�f�$!�;�`W\ O�gz�3�ӊ�B���� �R�U���`*�����c��������dR�ȿ��L�?�������k6@G�ED�(K@K� �f4�pF����Hv�)�H��ǘ�k�F�_�)'k�cyp�.?�c9nhh��ϟyf��Ϋ�}����緓�1��ftu$z3X�P��~�=`!E=�;F&�L�t��py$�� *� d�h��NJ<1i�[��;C����U)�?!���&���];:�N���(�D��ׁ�{�Ll���t�����������3&��ā8�v")��vA����[x�.��(��4g`����i��U�J����![���=����t�����65���Ķ�X���9�5& ZSq�ѷ�C�5#�6��loC�R���z���2��������t��$
�?O�Ӗ�|�����f�п��?1�(�o{�w� ��@�%E�"���Q�Ն���kB�
��KR<������iwA(��@a����&o{�͵�`s�?c���	��c��(��^��ch('�/�+Ĕ�wv��z��xf<��耯�;ĺ�(���U	��!���?�ص��Ϸ�T<��I7O�{a)�.r�-3@�PW�B���l��A�)(Ÿ�]�M���9Zx�Ș	�����>��������W6��ϕ������>����W��f��k�dr)�:�K�8�x����7�H$|��I��݊��������~1.�l`k���3��/�a��+�3������7�/{0 ���X��<�/A���\ny`�� M�Ȅ���ƒ�?�w��a�L"�d���3�!�}�
��_�x��'n�����^jwbZws ��k�@U������zs	E��"�)E�������ߟ�QX���0���\j���gFw6��j����$��_yg�Hq&=�y�ͦ�����H/?0�A���4��`���Kԅ�ƽ u�&;���e(58���� <ĭ_��­￥���ē�|FW�� kl�ˠ.�҃k;̊IM_҇#�L��zEԵ�VaQ�����*�c�����[��^|��|��=ӽ(�0���6�'�
�A~f���`���P��8\q����Z��^u����9p�K|<��&��c�;_�D�?�}0�n|����O�;�!&��"��]d%�ӥ�̚��w$�%�]X�%)�`�V)�w+��x�^���ܤ��*!l}�G��y��:(՟��3t0G;a*�r�PJ`z���K20 ����n�vf%�n)x�q/O�-�B,����S�����G_�MG���w��<�:�Q_�{!(�Lq�-��%5�C\��9F���V����l[�(��b���;�n��N/s��&W^S����|�$��m�So̥{&6OS�8��-��V���݌Yqֆ����J��,��o�+���	�.r��7��4zɾھ��_�>.s���og�נ���������%�`b{TX;� ��)	�Zq�X5�]�\���i��6���4�͵�_��{���[��\�gz������ǥRD���k&X�(����SH�,�H���-u����8��E�S)��C�1:�W�ٷb�G�W㖆:FH}@�P�6d�hK�ԛy�>�He/QRʀ�S �	;
zB�M^��qg�M�����w�c-�ۏ����^�����
P����Z���fT�9�e�� T�W)�J�{Vf-�{�mI mݢ����р�^ *E��Ԉ����w; ���0�~pgfzb�ho�G��s)[H֖1��@����V��aS�j㾬����[��T���2���t�'��P��#�͆�C���W�j1W�� �#X���6C\Z9��7���{k�Ϲ��9.�w+�Xyڣ��R�����\�N�"�9�>�֨���C`��E�������= &�O�Lgm�.��
�B.�*�LrP��*2��I�+�:�����H�(�{���<�pډ����"���ԙ��P���wP'��HJ"���LO�[++C��A�V�ţ/-d(ۼII1��C�]��0V�J�5�a;��&E© 8����U<�#R��4Ž��� r2P�d�
L
�~\���K3�1�uIn)����.u���<S^��ǓǺ�R�n%܉;��.�:233�&�9���s#�'��^C}��o��Թx�h�{U��Dh(�$�x�k��>�U�ʑ���Uq/��B$���T"u�/y p���#05��c;v47_�������NRG}���"���������1��c���PeM�[�.O�U��֯�ĽԿ+��"�d&8�GQg��I<C>hYh�p��L�?w��WGwUVV��Z�PP��P�\SA�����]�2_I2��4�e�]�8��L4�S�	C���R��}��3� 4�8�]��å���_�)��_��Wu+~n��s�̹v�%�]I�I�7��4�1L��:�;d���c���?
wD��� ��#����͹JhH��R�w%�a�0��]Wp���}Uԕ��	�SЙ�H��x�M�t��&��R�|�h__�?Hgt�OL�>]�:���ǂ�>6�_���J�/�zZ��m���E�=ъ��-n�Q[������5Ή0�^�Ag~���}�UG���^��M�������+5���G�WW��%koٸ���j�{�nV�t���vΦ�
4FC�~�)oh`W�m0��n���;C�P������)��Y'����k�=�w� y��I�������w�/��v����G��L�B�a
OA�C�#R�_���o������u���>�i�������!��*qy���XN>���U&	����p,.iz!�k;@�qr)�a"C(�\�%�[@�Co������{�����t���ٷ�5J�R`�%�%ٮ�����|�
�kIL�~����(h�	�B��ԧ�S�X���SY�d���NRL�>}������t�׭�!�;^$�,U�V���T(-�ʊ�+�]�PC!��2������'��Z3�w���������P��{����0Cs��wJ�Q��M9�<6��!�t$.'�ׄ�!�n:���}U�ML��G�*#�w�	��?��RRɡa�$%�\�|�RP�� �C��]�ч����MM���_k��m� �+�ͥ(���z���0m/���;ۆ��" (����q �,"�%�J��άw"�D�AK��@���_�g�P�sw"����ÿk\����멐�	�^��RƪYL[K_���*Z`�ESY,|�UD�	� 9e_����n�����&#�Y^f��D�.�j>Z*"�Ti h��r"�T6O����9����z�|��_�	xM%J�Lٸ�Ij	G����cN炏�b��s�ܑp,�P��b,sN*���\؉l����`(%IQ�tud��?�s'���w�2��1ћ
��R>Ш_��$:ߩڿ��}�}�A]uvi���L �vGb���X�]ik�r=��b:)��&�3�tU����*�DQW��,�@bp�����f'��;i���w���u��;q!�o+�5%�Q�c%��Q����Ĝ� ��[��l[�0�k���X�T�2Ws+S限0�ֲF�afV9����E$
ͽ�w��..t��׸������F�z�(̦C!��7���Z��2��e��j���I�Ӎ{�*�Y�.�BE�g�\����� >#��-��.�yi�Ѳ����	��CՔ���?��wX����F�0���Cq�NႴc�FI�W��+��҄{�>�dN �+BK�� ����`O�(kD����dd�E�0SO��q�6�k9��~����w�&h��P����Պ�늾Rd^�f��zu�3(�p�J5��r[OK�M@�H ����T� �]c{nml7��D�B�1�eౄb!�B��'�k���g���d�Qa&zk�ZRʵ��hIG
���e��M�#h�]Q�ɚU�݌��=���l +	KmY��@���`�=۶6��Zb�K�D�8�:��U	�μ}p���O_��`?t�gӸp:zKR)����+��ˆ�Di����5���M�Y>II�Y�.�{��� ,�Z����G�� �AɦgpJ��M�$��v�¨\��b�Z 2VO�"��d�� ݟ����Z��߅̠a��g�q1	˨S��!�l6�|/*y�Z��2F�k��ܜ�f�=��N�+-�,j{aWv�����V%(S��Q��]S
����!`V���8�`SO�hމ6�j'p�np�"���,eX�h\6�ڙz�X�𔛓���
Y����d���mh;�>C ��ٮfċ��Z��`&9����"V.������Ѿ���끛����>����=$J��
!IE(�v�^�|
R1�����(�g���H��Y�e	���)��.��D�!h ˟Q����kLI���������;��"����kk���-'����<�3D�N����j��Y�+��k9�+�� {�4Ӷ�(3�2��Φ�)5 N& j�ަ\�g� x��1K�,?"v���Uq.����W�����n2�������z+'j�`�W�e�d��T� {j����P�b-�ds�$��q�I�RI��lmW��r��FKyi�Տiw��vc)6a�s�'S�tZ��-���u��4ݫ�ue�L����C�^~n@fb7?^f��o!��*b��d�3�TĦ���,{E½�v���;��R�ld���G��qa2蝑Y6�t��(3}׷}����艟��8	�_"M�
?�ͅ)��c��e��;s��b����\��Gܑp:�T���9�JS9lgY�"�)�����.�Ƃ����(Ѻ%�[���(3���(� 1�E[���LAl�o����^Ə��gq�M�g���,%���x�p��H��i�bq1�#�|�	Q�`/N��f^RC�L+ u5�n����cqc��W���զC�c�41������K�w����ª�I�&���<G�,��b�"x�A�N�rW9�R��I�"2��Q�jk���ɒQʁ�*]�k����E���oKޛn�x�
{{*���ˠ�W���zS>�m}��	pP�K�}����{8�U����{ik�l	u�ѿ�����Aھ��/��H#O�˫�Tk�1��`�����;���{kJ��QG��pAy�Aq_�I��A`3��
h�6�O�h�E�����-%2�U \��0���xb
��۪�ߟ���o�v�U&1om�8)��������S� #Da�Ѳ\N�l�k�qɥ�I\��P�}�Z02pD��0�۸Ϡ��tpD�Z�ښ:�R�@_�a${gI'`�R�w��������K���3�w�{ �-Uر��x���F�w�>�\�K`��I�b���Sއ�H^2�"�\�w�U�@]�[�I���"2�E���J��ेS�H�ؖ._��6��F�I��G�����4$��)���[�J�/�޽��a�޲����v�>[T%|��� -�%^��Z�"�;�WL�VD�����^�Ȩ��r�@�8�#��X4&�����+KUI���xk	���Е����/�����c,:����*��� ������^�>�-�PJ������ ]n�%��!�>�i .���q2��ӍL����$�('Ǔ=t��3��Շ��Q��3
��Iq[%����{X����7�x.ҮV��$ژ�]�(��L�|��k�n�;�wu��w2REK ��b�ʝ����JZ*f���qWT\N�����ej~Qw-4"U��V�s�4c�4R��&�X�䫢��j#+?ǥ�wRf�^x�^L;ba�Ke����)�v�P��=w�@{T�9�?kD=����U!�ɷ����}�R�=�6��b�'�܅�=?JHŋ��E�KJ&?�G�����|v���i;�'A� /�r`IK�R4'���à�Z'�{����!<ի�<+��߱�����]��|m��ĉ��IN٫�ܜ/דH�튔��M&|�{|���j�=��n���D��Ӵ�d�6�F:���plL�-A$���eWw�`)�����PKM�>����i ;V�r!ڗWK�c%@�~g����l����nb*Nʗ�vQ$�=�S9Q�;�r<.,V(JO�������m\\]}w7�,�q�&8l��&��T�c��6'��V�~�댪?�%���X��0d�����=�};��ts>@o�DA��֟g}ݍ�Ǐ�p�uuuE3Q�N���)�n�lN���I��e1?Z�����bB���J��Q�z�CA�<w�^Vm*ϐ	�?8��7f���c��	��;����뺅w츉k�Nb����~�2�Դ��ؾ���z�F��jT��'��ϺWD��y��G���� �D3J��!< ��`�$%9����.f�bO}�B`R�&1�߳��D$f��	��jvɰ醟�5�p�lJ6F5��%�[5�p�D+�.�s�(��cWVu$;�&�W3��A(�� ն�1��7uf��kG6�Q�����a�d��v+a����F��8%(U������f�`ߧ&qc�TOn/�����Ks]�tY�ˏ�S��ۖ�l�k:���3~Z������g�D(5T	�������f�������i�lM�F<=���)�^6�i��#׮��<ܰ��8v���ޕA�%$�~���;��x��ES{�n]j�L����@(
3�j��$�`,�!��kB
B��N=̥c�.�&������K�Z��3�B�������h�����w�X����ct[;=�Q;K��vz^E���ul��{n�a�126F5����k�S��*���NL&�:�N�Iw.��O����'xٲ�O��'0�?y��*��3��
;�&�̵9���3�yaB^U�QvU"q����f�U�x���B���vjw���8톖�eF?Mʨ���zǁ96��S��]]��{)�Y�	�`,��I{R|驤"�IŽ�+J��%����@bf|Ɋ�e���-�OI�a�����|W0�ˁS��N'����/�}��W%�㲹\C��`��~��O�wNLw"�Cq��W���$��q�D��n9ra��8<F1�	�͸%3�e:YpG�E{ ����4�tΞFS���/�ӗ��/�=��>��L�&�Q3����U���8�� ��:,�i�z"��ű��L��>6��{?zb�&�����e������8#�V��k�(;��7��uvv�Q�ѝ�:�<�v\�O$�S�`G�z*0M�2ՂG�L��zf0�S.WdgH�:���%sZ���
q�-�@w���?�N��/�NT��p����6�m�X3�oz�NИ޾c�.���H�]�GSa�JyL�d�7>~����Y��X�H{{��1tdV�G���
�͢~�&!	z&lr
�P��:���3Zf ���6]�Iu��9�\$˃N�ML{�W�0G K6�*l	�0V���k�# ��Ro'6ӬO�D�ʹ��i��@=��`_?��Ȇ�G�������H�H�	u��kD����s.�K�B�$�?-�\����mˀ.(~K�fX��ƤL_(�4v�hg��1m��c� �ߖX�:'}�!q�m'��m����N��;+�Aى"
=Π}Ʌ���z�0��ۥ��uGnn�y�1;���l�2���������}&pq�*�nP�Xx�M���JF���p��&'h& �k��P��.����L�ئYU!R�%&��HB]��>2S�������/�B��W��)��	�T�7PoqV�+�̰}�����@��u�#c��|� {��ά��z��'7�t'�r���)^��Ź�D�넩���:�Tb[���%�sd;�0m�t��.8l�yP�����V�A����nn�x�xL�K�] �*h��ss �S���N�&�k�.=0��QL�v��{LTKen�D���z��42=l�������{B�
���'U�D�%�$��r���T�k����7z�^@�#�����{��Q�8�zX�K��8r��ܺ��Fd:"����ս�d����f{��o��.�Z����X@WX���������m��~m�"=Bc,I��C�7]%��~���`W�xc���/�R��t��צ���^�H)��]���~����$�GO����7o���n��l"=��n��F~x���~�l�߯��#�y��?"EAN���	p��4ͺNS1Y�O���n�Mf��WA�q����S���m�П.6�X���kXW�d�3�9��2e����!��x�g��'�t���`ޱ����=:�v��Eo֘���.�e��zFxp�����G�L�6��b�iޑ�$��'jCl��qy)浻9Q�bB���=d��Z/�xd���M�Z����ڋ0���4Y���I��zoxJAix@}�@}����qLTʻ���Ý2ю��6���d���PfmT����PE��\L!>r�Vȝ�x�I&bNo	�����.�@u�����	��c; l~�&��^�{�u��x��.<�JU��񺔨.a��M%���*1��]��w�F#v },�$iO��\�o7㾦A2����D�i�_ĕo0�M��x�yG5��m)#����B�:�j��ђ�D�m���t��O�,#h:�,]@�F�����<�̿�Dϒ��#���8�6�6v��� �<cE��?<<ܘQت�G7���5�N���S_���}1��M�;�� ��#�u�b��&b����p샣gqa�m)6�^�;�nA��;��	���r�u궰�7��&g`���_7w�����}Lc{W�������o�ԅxX��I+���^���'�f��Qԝ4�h"{T�n� ���J��W�]���m��M���	�݅W9<�	�x������e�h6���vg�Pk(D�Ay,t�U=ܨ�D3��7�n��Y��ELgأ����,��Է��E�Np)r|*��D1CӝF"�i��[a��it=ϋ�YaFe}l�I8�Qe)�����[ �}}�*C)��Z����8~���(]{`����ng�nU�F��4��a�����C�՚}{��Q'2ƕ\֙[Խ�b�5��Q���fϨoۃYY3G`�+�lX���O��[9t?��7��)�<VɅ8�m0��Qg�mJ������7/�u/ɵL�XƂ��F���C�N����[d��j���"��ӫ��Sީ�n'~�Y֍El�v B#̨���␱4;n���@<^N�̡������fc�8��i�����`��O��7�߼���ٰ0&�i�����|�1\eE�������%RBu��i�=d�\'�SO�b*&���,ђ�IRq!�u$��T����F��e�f���_�R޸Kٖ�I���/lD��7�|z���@^�����?��G�Z��2�b�X;��T�
A�M�[�z�|��"�5=��L�v+ȧyXkTM8�ݲ���UbmO�]�x����Ky�5!.�+����!�k�5��u[���T���� )�8fA�g��#�+J4���)���fd�]��#NS�Ŭ�x5@b8��s�FF��<xif��-�"�����y��Aǵ�����k+[]���B_��Z5i��9����$��؏�t�g��
�U#E0Le"����,�V���au��*.�b�zΚ	0l;ͱc�����Yd$#d*�! �KII�\\��q)�{����?ݛ��=�M�3�X���'�of��=eط�9F�4�h�UoPڣ��^��'6��ਯw��R�8c���6��8-����`�I~۞Yd��)_Rf�$&��8���Ae�y���yM�N���1�O)':Җv�4f�vu;�l8����E���:&���|LUEU&*KQ�6�F��C�v�e����6�}ў1]3�����S�����]��]�x4�_�����gpR]�� �_�^И����o$�]oN믻q���u���*KF}�QG���=�b�Y������|�"�KZ��p�������	�i�k�u�	|L�Y(.�1U«yWS<(윪�b��L�-�FeW�k��Z��<���G��7܄�nvds�l�Y�����c��͋/(���p>���?���� k"��a�݄zA�����9A.��YW,��
;+�WE�����!d�����G}��Jn��-l�*d���u�1��X6�b�q���F���%�҃����J"L��Vy(��kJ�$��t,Yl{-~���G6N��il�i��ݱ�,e{����9��+W�a��7�;q�5nT���zM�p+��?�`p�4vi3j���ZB�����^����*n �/�p�u��XT��q��,F�
�3�ci�F��s�i���&����<���a~1�:�c狘�Y�v&ԗ��uv�*���F�{���︀i�Y�V�h�<"��4���B��l9��ا��L�+ͷ�����q��6\����"=ioX;[O_ΰ�L~Nտ)Iw������J�{��}����umgg/VV��<�=&�ʾ�����GXF �ޮ�Ϩ�z�9���<���A�4�@�[Q8,�$��V�1�Ɣ@,Kq=��Dұ�eN�=k�L���dwsm|�`#�n&�E��_�Z��Ͼ����W��7\��*�̀�i��~�1s[�#Xʞ�H��	h4�Q��S4�)��ݰh<Lw��ҷ��I����uC�e���m��"�s[�wBdvF�s�^$�p�f�B�Q�ؒ)}��`)I�{/E3دp�i���K?��<�P[C�HBO)�Qг�<�k�۩�h�J�fe�2��%�t��ʁ�$�N�`�%�}�Y���=����	;r�-,��1{�=��ذ�r<�%A@$)�!#+XHz9�.Ω!\�Ow}И��J;+[�Cq,1ͳ=.����s���c�V%����Z�7�ݕ4.��q1����{Ñ,/p."Y0~x�I~_�MY��t�������3����,g2Y���&�d�wE�Ȩ�3�2O_���+����|�;=щ
Z~m�C`+MJ*;x��ZQ��,&_��	��2|U�^v��GbZ|�D��H�ۧ|
�}���P��� p=��5�-�"��Xn��	����Y����V'c�i.�6��>��ߏK�;��_�N�M3���K���kvp�Gjw���a�����c��Ƙ��#x�p�XT�b��ZV��V0�)6d}�dj4��l7�����ppz���)Eݞ�}q?�Z�8��h8k�o��JN�Y!��x��i̇�P�ބu`�w��B!ό���a�a�^���٭�ٷ:�M�1�I��<�R��%��]�	��A-H���§<l���6�	RFc�"�ޘ�(eb�7��G"��$a�N��H7���gt�bڀS�����11�t6�������=3�Q[��&/�\��u�3�~ށ���u�v��Z-{>70�+{#jL��k�u�I,HIǊ�4��(owsy���
�[��,T��B8 ]7�dS)���V����%`����9԰����x���e79.�6�T?.)�6�8:j�[CbH&�ݒu[&TɃe�nǁ#Ǐl�c�彺�4��5�����5L�H�\��zyJzg:�M?4�5�`E:����׉�Q����"\�@�旵�4��$�3���؛�y��`�%��,%y�Yw�ej��_��[��t�Ψ����������y�2�2�7�l�y`a�a"�1�60%�8���ͩL��Ln{��<w:��4'���t���Q��ۈ��'��u;Z��0)�i,���s�
��X��|	���،DB[��q�U�+Q��?����k�!�)-K�ѫ5luQ���m�c4q��M�nb�r�>��E3�^����-0��싁p��c;uBeh�#K�������:ك�T�"�`��i9L��-F5��Z����V�ї����`�{�����x	qo���_�'������1v�1��}���1tJ�?����-F��L�����]J4��
~=�m�T����)�m��r2�Q��)o�n�ǼE�D��t2�	�}V�0�n�ۼ�WRd$}y[`����}��,$��z':��+S~�-����m���.�Ú�g�:,�����ZS��� iٰ��Ѽg�Nb1D:��`�Y���=��PY��C��V��A�=��c�������N�}��n�\"T�S����C��_�C)q�u���鎎�+C\��W;z���v!�9�e���Oٌ:fJ�`;�V�2]�"�=W*�J�AM.<�KŃ�8f�ǳ�X ���	�� D
ǖ�*����v+��e�5]���tW�"
���/��CO��I��T��x���Q�������]�Y�0fw���7�}�qp�a�U�ޒ�m0�Q�y�𖕍2�Є�*��3�<��:�ρH�-�v�?n��s��k��X�oI4�=��%>��P+�1���`�O ���ưS���K�	Q�3�u`�74�����kFr���L���i
W+�`��{,v9���*{���Y������XP�]s���t$�G|qv�g>�M2ea��ZJd����R����?*�y������W�+CbܥG�'-�%�my2��z|C]q5u�H�,3�ߗ�x#(���E��(<�~��hq��Y��3���N@�p}�02A���H�=\ 6������ZF+�K���D֜����X�Tj���z�������+S!?QL[���#���� ����b�k��z�o#Þ�Ͳ��.��9����6N~ �=b�żi�*A�-Iމ;�A`rK�8=�S�
if�ř�
�g���o�zIe]d`{H�/Yh!�6>�Mm���C!Q�^] =�N��o?�0�^Z��\�L��46�7�5�aN݄;�<i\��-�&�s�H.��PMݩ�R#��w��K{� Fk>�k,�t�?0���o�2EK%&Uɜ+(dv���>Q�e��ic�"q�u��wk':@�[C!������8�-2�h� V��Āo�H�/�3j"�ϭ`�����2��B��Vd;�����{��nk��� DIX(T�M��px���X"��n�r5&?K���%�^zޤ�!�o"���08��Kgv\��dE���Yc��r/s����������S�ͥ�k���y�;/�W�(#�P}d��^x ���*pJڋ��e$j�5�:JXl���)�[8.�-�DӂRI�)z��k[<8�a?���\��umh6�	��*��/�`d2�7n�ܰn�$�5qgv]3���'��@{ ;�{�H2�^"\2A��<m0B�_�KM�'r<����.Ou��"弋���d������s4�hv�%E�hV�L%c����P��i,��V�a��o:Q�wU�D�W\ֳ�N�� ��7�����x�f�kΑqC$�Tbh����,ϰ���pB(�h�~��}��m��<p=��U|��ZG=��o}4�'�#�4Ͱ&f���$v`�����c��ݪ2����	:����n�/��/1��(-��Z�8���ۓ��]��6�Å`^��ԕ��U�v���+��\��tf��fm���K�7��\�:fh_�=��O�����HZ�Y[B��kHj�Ȕ|{h���=�'�B\LUm�V����ybbZ�Q���.����`�M���|a;?f���)�-�� Ց�2tÞ쎁�Ic.�Ph����p�B�ք;f|�Ң�sT̃�
���ڗ@֍�h���L���Ș�T�/鮺��Ip�5y��C�^�V�����!�|bf�*Q�:Ad�t�������\�N�FVZ��b�aM�qf]�2����M�ѮLΪm���V/�f08�)���p]�Da���vgP7�����\��el�d i��Jmv�����q'�\J�j�:D��{���~k��_���΃C�P������q�e�F���sǏo���|U��_cظ�%��l�0�`�v)m^/��/1���$Xp�Y���d�$���X�-ͦ�w̱�p15<�9��!�`�����(�ɹ��tQ�#�� }�Kƺ���F'�(��=ُ�x�S
��!Q���z��`�d�f�^�S�7��m4����d�0m���d��#�tZm�f�-XsK���aUM����_9�cG�D�6b��]M`��T�io����"SS��=a����;Spjyg�쥪����=�:lǬ�Dqgs�I�=��k��;6���%x�##D�g/`_���%��l:�7��ѱ3}��1���c8��j�X$�i�ۄ>��@:���e6�q�R̦i�+Aͧ3��0#k���mS�M��!얝��� �ҧ]�ELW��N,���`�����Gq�o�l�?��Kw�P�Z��gd2F�W�t�n�̶[6�7Z?!���.��b$ �)��t�����׋�ˤ�As^V�ե�Ԟn�.��'������1��.�hjLSf#X����Y��h�+*�cZՅ���&���+�e���4|�2�������?�mX-��a?΋��m���xıJ��+ș�86��>���X����P�a6�훆�e�鄐1��a{��Ur�X�{�ki��N��Pb�º���3s�H[Й%��D;�i^ݬ1x�6��q���۷Uy� =HbM�Îø6��|)�{ټ��E��!bz�� �?6���6����������R��Ѣ�v�}�(��2��Heg_�uMfAj���1l��c��^��ڀ��6��u��
�3�$� JB�mVVI� �@ �Ac>�µ��)\��(�(1��j�Ec��5�����{t��D)��m�vm���{�g\�a���?�'�n����¤^<�W̟�pR(P���u7�c�4V�o]ch���ԡ;F*-����.���-8q�=�^�k�P��C��y�=x?��HO�y�ӈL��Ic���G{p���j	�L�&e;^Y��@P%5�v�7�~����i������P%�2Ɯ���~Z�I��EQZ���{�n?~����za�t����]�Ff�ٻ�ilj%;��r��)U�1P^�ٱ�)Y`����vaա�'�a\������
L��V^���+�ȍ�!��NE�B�R��D?��2]E	�"$�U��
B ��=�J�~��ԦG^x����յ�8�H���Z�x7獍�E�7�=z�T4��w�T�K�0�//�
��pBE��G��q�"3�c�@��C���de]Aat�����mí�� 1��4DF͋���KA?�r	�K���� 9.��~aT+��n���jC;���o+sh�7��`�eI^�u�����fq2=߿�_OCv������~Xۯİ�1�a��0�����ڂ�@:��u��5�Fosfg��Ng�^M�i��6p�^�φ-YŐ~ʕ�)�N�.�S��A���xh|p�O���ipL�@�C��L��i3C��"퉰��adoڸ�Z��\�*�j��z� ��6`���̌564�t����oohXn1*~�)d~X��lj�N�Û�D��!��ciP���Yf���1o�*��ys�6�mM�v\-�'�Г^F8�g�1���X����|�[{cpy���������j5��W�eⷵ��D������6������;`BI~�V~J�l{���#�o�����m�g���v����EfX�+����0E~�����M>���o8�O��:�f�Y�Z�.�����`�^��k�I9�olFă�Tٯm���e�sd��D\��g�|�F5��g�>���.ֲd��c�=硅�hx���~k��-"������T�;�����7��j�Y{�O% |a�ISx�s����#��#�����w����m���n��kyd.��&�G�kdx��ѝ�I�����p�o1fn2��~��sn.<�',�

�g���#�7¥�Hd�N���\����h<8p�9��9s�wo�� ��_~}����Sx�����(�&'��t1�iC��?rw��V�ͽ�=��['~����v��g>�!�59p~��ܰ���}���q��}daq8@�#��̌1p���o��'���/���E@x��T������o&S\��*/�+�^D}�/�ZL��sK�b�Q�)D�_:w�z�@<���|�r~��ʩ3[��S����[[���H�K�RC[�ͭ�v�ƍ�{m��h�����w�xD�7D�`�������8�{�fӘc���͛{]�cv=j9[Ke����@�k7j"p<̭��6��'ɱ����J��_wx�g�̂!� �x�,�x����QՕE��?.@��^]���ٚ�.�xu5\�c�'�ǯ�ۗ�j���~���������掘�ԏAн)�@�9�;���+/�����B��[C7�I��DT{?�ܯ���ݒ�v
��k��Ϗ���m���׭�0�=�d�������lb]:ɵ�
'���h�!��zu�I��)�d��y%QG���� XH�Vqm��P�n'��E�8h;�LM͝3�ϡ���߽{w{Mu��O������w�|�ؕ�w_�{g||Pմ���x2튢��G�><=85�+�������m뭉ξ�PHT�˗��x��ۻ��q��w����Xw��c�ñu��, �wl�v���k�@{������e�R�7m�6t�zCr��"����a�4Pj<�.8��Ɓ�
�XJ���δ9۰X}�42�Y�S�j��U������r�n͹�y����f��3g�n9w����N��{��z��3w��1>(��֍�'W�U33nw�n�8��Ep�4Lmz䫿}�sd{3���@�?
F$��`Ǎ�0�ި�p��h�u`h�c����u`�mol�����(���u	G@j���Z(���`v�A�YW&��؃�n.�����R~���hsj�S�.]�~jKu��$�<z��ʖ��l�9w�җ_^��se;�~����N��JƓ��D���l��K��Ŗ>M�l�ɧ{)�٫ȷ��|��~�fd(��.ԭ? .�����ٺûfg����1ƶ��
~��o���:����B,��v�9�Q�p�O a_��<�=�g>����l{n&�g�ItO��V\��)��}�~p��-�oJL����s[N���r�Ԗs���P�B��.�9[��.H�W�X���)�(��	a���
���3�e?43�hۏ�Z׍l�E��v��� �o\[�`� �7�pt�t6��Q�a�if�V�$#`qZ��ڂ��͖J�\���&�2U;��F�TS"V�c\,2�`<�Ծ/����n5h��6���һ�^͹��K�w��3����rj��j��+�/������*=K�.�~���q�K�󞉫v�^�u�ڞ6p�������݇�f���:;�`w�>|c�7v_; :��V��(uy�`l��
�n&��Jg:�9����w����h�e��/V����ap0t_����"*%��6��ԋھ��N��2~rP�9{�̾}��a�W��Y���/�m���_>��J� s0.���:=C�e�$Eda�v�i:�������t�.�=��oY�\Xt��(h���u�BF��}�an ����6�;�����F�
+%yײ�tӔ�4�@���|BM�W*�(�0
���rj�g�h�<�i����ɪ����5��f/z�N�_�{���Հ����N}�� ;�HOuu���_�;���_�ˬ����.���X�L����H�GZ�VF��։���-<e��N_]�%|���*��]�R� ������n8f{\���#��Y�+Ү��Tw�"�ł{"/��W#��ߚ�[2�����h�nf�1?�,24��L�ԳW@A���1~�.~s�җ/�^}���\�r��������Ů�*6��:3 ��H���{�"����nz��������L�I��
�ɔ��y �%��.�B�u׮��{���Y�~v���# �#Z���܇�N���,3�3TB8�B0�� wk�1�R�H��*�~Z�(Cح9��"�.��~�F�g�4VW_:�r�z�)��[�'�Ξ~
f�q���]��i�ͩqqw$�u:�س����}��>��:'6�֏���Xg��";r��k� �av�d��9<0�o�� �.���Y��ǰ�C��q�U�V�7jl7Co��X_P�����ө���'��1�.)T㉞n�l�XMd\��;�6�lu���H�;�^�o9u�`N��1�;KOl�ģ/�Y�p���;�px�q�_}�9�y�®UkLz������7�V��k��=�V
;&x�@�^�oo_�~����h �4l=0�>�j4��خþ"۵�_��hbx�l�G�j��%Kz�#�^�ȸ�{5K�݁����+W��=}���ol?��Җ��s�N�Rs��s�:�C�<{�d$��R�g��h���>훘8��NC�DڛNʲ�N{���~�vܗ�/�M<�q�$��µ��`l]n�9U_�f�1���v�aw	��4�Pʣc77�Х�*�*2�*�%�O��>��%@ƩSgN�T�W_�wa�EwsC���yRv��N���,x�I���/�j����|�G�d@��i��;���%�7\�0p�u7n2؁���7.��w�1���8��ՑYǺ��>00�h[f�K�%���Y�vBϏ�ۼEd�@����	�80q�a�L�� ���0��0����Q�x���;�/��l�s婳�{��۷_��{��=Wgޥ����Vx�<GDq&�bO���}�}��Г��ٌl��C��1owkq��6�B4�uƔ��=�����g]� ��,.w,��;�������e��ИM�h�J�w뢩&��3�����HT��$
<�qԼ��R�{���D�~\�_���a�ڌ���7{�@o�K�Z�� 3~_8�"��=Ty���}��.�ڤ��{+2UQ{����BFb��ߣۮ��w��5��c펑��1@������t.��_�j�0B����%�*�I�ymJ�}�H��UNe[EF-Gdp"d�j h/r��5J�C�-x�ŕk"c e���f%�x�7�$\츀�7���3J2�c�%n������ <�W�E��!��hx��Bk��z�u	��T��E��ޝg�N�-��QTP���Q�Iܖ��E�1^f�'tvſm�ui����V�r������]���O����y�k5�3�;��/��C"� ;�9]d��g���w�;u5B�&i�q���Xf��Í���a3�K�ξ���|��'@b|����G��=Z�"�j��"C��,wE傸8k3�3V-ĝzS͗�qp�΃R������缁$G x�`���n�}a1��m.f�*^�v]2R�a��e�Ah��"L�}=B���t5�+J��EKK�2�a{���v�1�3<#�vz$MƀhuDZ��
F�~"C���%V��b_�0a(q��l0=�x�n���޶�N����Z��«x�e{s�~�u�Aځb���`�s>M��	�1��ͽ����a�g�����پ�W�`e%���)�:QP`h^������_��
F�>"�~�GY����E����P��y����ڽT�3V#�a�/,��$��S����/�v�pEP�9o07�ڮOy&�g̍��㖒�Fm�U��Rd_���M3��	��Pqv�`�,�TUK%�F�Pd�.*ZI/4aO���F�R��$�u��w���"�{Ӽϊ����v�&�dn�Ϛ؞���>B�?��[��W�~��ȲV��fS�w���lN�8�\Y	w}F��SB������l�L撤7S[���K���6�Re�TU�:`��Dg
4ohzQ�,���Hr1��z+�v������kf�������|� ����m�>�e~Tw�-����N��ƱMt9���H����7�7.�-S�^��T�qx��r�	{`����_>�@m��a��]�c�AZ��D�/)a�AV�99
�������I�fЕ�}����y����'�&qݦlW��v�WQ��O>�]��B��d �����qy	�B�ǛNhd�-h�ݡ�7Sww��2|� u��q��n�Ý��6�e����]��!�Z^��^�w���#�켇��^e�I�=V72.}sa���z�c�E99>�:>�잇��!A�����i�ho�E���_+��b8�s��&�����z욶�NO\�a�9���>����0�k�Nwoo�u��u�l�@������?0P�bVG�z��F��[6�2x#��v`��o��Rq������'C��}��������ʚ+W��ܫǫk�l�R]yr�Q�US]=?X�F�̌��?W��4i���rO�)�9����įJx�U%������k��Q�3ė���=��y#���%9�5y��tݍ7֍�ήۺ��܍uG݁�׮� 7G��7����w����[�G,eaIy`�w�P�}��.�Qi�dx�T�������R�ҝ�o��~�̩�X����3w�^y��-g_>wV��q��vw��z��sg��5��l5O�|�%opJ���oxI�,r����Z�>��,=��n^���릍	���7�P�Yf�c�����l�����#����^�vm���u�w_����5��p��v�c̒���r�5k����,���^�����3b�kd(��b�W��r������>u�ܖ�gN�:u���+�.�|z�)���sW���;O�9�k\ĦYɳ�Ճ%������{rx%V[��B�QdpQoJ�>��������$��8�k|���{]ݺ�k��a����:�7\���X�1⨻q��@�Ed6�:�W׌;��h�
>F�X��@d
�7gd��-��<;�{�}��� �\����ӗ���w��K�|z{͹�}��w������K��[S=H�����lW8�����i�PG��3ط�OX�������i{����Z�V�T��Rгw;���p[���{`= �uv�|��+p��_�0wx�A����bl���$_y����i�a6.N�YT�g�Ȭ����������\��}O]y���jν���w�⧶�\����W�|��+�����������r���m�6��bξ8��iͫ߯������D����e\�q?(���ޏ��sP��9f쾰`*ߨ��[���`�s�nd�:��.R�������c��P�6�M�g���X��{�ԑʱ�r

gD�`lK�B�_V)g�;m��:�I]]oƒ��a��	�<��b�v�(
H�N�Cz;I�J�?��u}>�sN���۸O��"��y����/��^���]�j9��5��E��)%Y��A�%�]�
�Wcz�'�X������^i��z��5�g��l�B(C�m��Ń��^v�N�#�!�������9�]������;��ƒz,�#��Y�l;�Omz�nߊ�V#�E���G�w�֮��@�̙�����&'G�ǰ��h�������w���ri�""��3�`����QRԀw.�H�e� �~�=fk�l_
/��7dnY� �M�X�_�S<T��Ex�1Iˇ�`cɩ�p���y{���a���L��6�6����7�,��\�Ns���������Y�	QK���t��Ϛ�)?��hҀg�Lɥ^ꀕռ�Ǡ�DfJD�o��Ngmm_, ��o��Eο�"`_�̨��ť`���^$��ˋ� ��0)�դR�1�z��R��"��ɨ֢��=Js䟡�&���O��^1k��W�����47-۴,;�d֙�$<uV'�e�~'ؕ8sٖ��|Z�Ɋ�����;�I�ɀ���ߴ�n۶W@�c�s��o��le/�RWW�
�?����3F3�<��}q�}�Mo �O#�!{"#�i���^�G�\�	g$½�}�ؑ��8^�`�`�[=�z��
�����`oǂ�1�#��<�w"<BeM��f�h�"�����)}!'�@��4��u�����,��_���~[͋�,mj�VW���`g"�N�_̄���NUa3n?��\dp�8�X��j���'�#�@b�+�\�	-�Yk�.x#��'��o��Ȭֱ#��s���=���̦��;ZOOƱ��U�O*�f�����~�5�ͣ��!2��"��1*�b?�)�> ���ƚf���1���������z_�v����^b;�n���.�?������~#���7����:��J�tp5S-4� �� 焹\ ��&�},��������@Q�
��OnbG�IK&�����t�����SMx0���W,3Tdg��Im��rY"��+��'�Iq4W����IY��R��_ʶ��������A���,#}!��tا�7���6I��9ۗ�/�O�n	؎�_KKK��nH;���n����`���N�"l�Y] ����:R�$�"� v,^@l�T��(2��Ik"�g�0/Cd�oI��J�x����.�����:8J1�Chɀ�n���+����W8�so��:ZEy�l�ϚaO�ι8<."�f�%��SvQ���h��5����Y�^T�~z���bs��
��="��Ad�V, �ؾ����N�K�͎!r�e>�4cw����F���#��0��+[���m�������s	v����>�SAg;��2=�S���*lJ�JvvZм�����K��#۵����7��p��/�ꎬ9yrN�3�k��wM�F�V�X��
�ŝq��}daG��<=�&�89�%��D�_RSh���JD�`�&Ý������z8�����	��b��ee�x�32�?���[oZ2�v�������[p��8��F{�׮���O_o8�`?,�����#՞������2G����F|E�1BP���^����#GN.�x;��G���J73�гRۧ2%{w"��F؃ �q�ݱ�:�x��/6��EG/lG�"��{��
`�����M�CY���uZ�� �����p���e�S?}o#F����b���,�p�Ժ���5��ճ�P(l֦՛�7�A�}�j��D��߄�^��I�9܋��؞�.*�GTQ5���R"��<���Qp~g���n�ܦ�zmM/�2�	���^;u ~3 )F��98�`��Xmp�c�I�mN%�y_�#���70إ���iODԗ����"._��ƿ6��XӺ�L�ɓ'����ذ�y����'ל��݅�N�"8����f��	����"��.)2�d28?������.��m�`<���+`��>[JNjy�K� ��%>�8fAdX�{zر�/�?Y
l?ц���TM~j6��^_�nl���/ _)A-o�Y�����Xs��mZ�cu7x��O�MY=�	&63�T�]����J!M�TE$N��o�_d����ɋ��co������/��_�����Gl����//��ߵ+f{}��&D��o�Ր���0q�[��i�K {`ڠ`�:��S�q���jw$�lvEPo"|�.WQ��N��Mz���lo_��+C}R�LW��}��#���;�L�˥E��`�����[�[VG(X,��b��������<}4�l�Z�4-�~�spy��r)��T&������|��[_G�O�y�L���l�Wk4jK�v���twuUb��L3�1��O:�_r�᫒���x�%ug���+G�~	)�)�!�P`�!si��H����=f���|ì����aV��/&kC�Ά;L����������i��4]��?�`_��	*po+�̸д���PQ�Ȃ3dʰ��]��n0
����G�%N�)�5�'"���t�Pu���f�V>p��ӯ�翆�J�*�\���"�C6��v�9]�Og�O8<�}�p�/�w8�I,��/�!+4[I��%�h(�%i��o췃�"�qU�=1��&�q�%#�d��`-�)�ͷ��Ŋ1���a24�W̚��O�hX����iuu����ӋLjZ�Aq�:}:�;ԙ!�v���'���'����%�.G�R��l�Z�S?|�>�����%���C	Z��r��ras�X��+F\N��7��M��Y���.�B�����8���L�)i3�B�z����|��˖m2�%���[dXQL2i��L��;ܝn��_�X����,5�P!�~���N�|T��Ё¾gZ�y�����ON`�F1���jnZt%��D�qw�v�g3O�L�ӝ�:��1��� ~ҩk���*�4��5���wVS˷�|���v%5������׋#���>�IvNy"}�<�=��N��pP��,��Aj@u��D����ġ�<�'��<��M��jΩ�L���ܾ��͢c����P ug�|>NY�h�G�l'�O���>��x��4e�� �����DF� \<�g��&��@ �$�;�1�W��/<�p���g�)�%eըC�e�p�C��l !��#��OfA��ֲ<U۵��ͦ��d݅%�R�H�k�;{t�f+��2��2!��N�:[�
���O_;�)c��R"��!2|Vx0< ��H?әR�4���m1�'�a����H����T��T����PqzR`��+���o����y~މ�66�
)�ŲT�c�(��!w�.����{#L�ɜ1u0u�Y��2�N_���^�'�K���Vv|�P�?��Ȟ��v�Q٧�2\cPf:u�mntR>�-�:>�[��Ȝ�ye � �1(C���ɔ��/O�h��?�=��� �M���t��z�ۋ\�H�e��K2�<��5c]��О��Nm���.3z?AN+FI�9� �ۇL��/2<[�Ɏ�?Ei��g��n7SO�N�OZ�
оTD�	w6����D����P߫7��K��މyˋk	��<88Ņ�cgv�#���n��k� �qU��g�����o��Q��q's�(���*��"���u ��@6Р1Lf��ܘх���a�Ai��x1|�ۏ!1����ݯi4�'�Bai�1㏛���<��`�C���̹x��L�9���w_��4=�1�#��X���?����D�iӉ:�JKʎ���ˇTc��e���p�&�f���\?R9���ܜ�d\��n�Xʖ����o�s8�������Ǉ��Sb;Qp話e�����~��/�S5�f`�&nB�0��qW�����d2q7Vu�g����2M%��(��0΁|5&���;����r�]��s"��rjN���#鸇�d�W_,�T�g��~KP�>��]M��L)1^�a7�D�}��'~J�W �U�V�ZUD8Cj����l�q�f�DL;��>��i�=w.9�(���:�!��L`hh��eDv��R�)2z�p�֘�#խ#�a������K�6wφ=�lɤ�^�c��zm�a2lS��w�vs�~
�~�/��Iy�/ա�e�A�Q�
ܩ�����U�T�;MM�{���tƛU-�$�{����ȡ���˷Ӊ����W$2�� ��0�a��θ�읝���	s�����ۆ�bI�x��ZU��ڞ$v���7�h���񩟞����68S�p���ʎ3^��;sf����$�'8ac�yw�S7ܩ��{�z����2���T�a�K��& O�v�|E"C�(1��e�3|%��;��}�7�-���6���CN��ƻK)IMUb� iN51�.����K�;��3eL47�>Q��/ qgA�FF�q'o�{�ۍ#�k��P��F)E͇j�����UH�_C5θb�����	�.���7�]��ǭ�ń;'���z�o�3�ߝ�\��N��� |%�-�����X���_}�'��.gy��n�{��k_6$v0y)�/`rb�$u���b��i�{W�%�T���%��cJ�0���,q��o���D��nc���󹾻��d��n᜚���ے��(����R8 ��3�<lǖ:Q3W�~����@R����U����ѧ\ڑ�Ɉޠ��qH�v�s�i=s3
7"�t6���{�뉫���0��DiG�Uv�f��/-2��Իrx�L_:��|�2e�(��v��=M��C����	,J	uf9����Zh^ܹv������z�����)�!6��8��##�0�x<R��d��}���;`��2��'�8ޖ��V3ԫ���*�U�Y���7�L'2����i�~��ԝ�ʄܭs݂�o!�)æJ�bn�aS8T��%����o�kjA��g�{+��;�~<S�_M#g٢ڈ��L�YK�d\h���<��]�9����M�^m��acΚ��#��R�s��~ф%����n4���Gw��t�
��Y�zOiE�ǹ6���Gaܮ���z��X�����1���^_�y����Qs���	�U�5�W��G�0.��)�N�:�9�'��3���JJ��h�Zg�`;#;L��ھ��ً9��6Sd��4�!���\���d���HͰ�	v�1{6l���U����7L�*��Qю������d�¾��?�=���Іgj����/!�McX�TĢh6�����tq�1��ɮ�gĴߜt/��2�D�[}YH�ER���"��V�iEF��1���,3�N��{:�1��nj`o���K�M�1��:T�H��Y��g��Ul�k��
�]��Eu�T�G�E�c���ZQ�dw��D�T�]s���ǝ|���TK�Dw��Qn�Ȇ���KX�܏���?aWL�{/-2��-��ÂGq�Pw��lϰ���^뉑CC�v��w2�p
'p _���fI;���?�ނ���ݮ"�~/pa}aA��F���5��>F� �x�GeٝF�=;Ƌ�р/�Fs�i�dZ�C���4�I�K�ſ$���,�?z�n4f]�{�w���ٳ���G�2�b�������t���qF&�k}�{�a>�PB�΀����7��ٽ`�e�"�$WՉn<D���v��������cE�Ik�zT��!�K�u�D��_��"�:���Ӕa�Gf"f�s�1f��=��|��}v,�w�����_i@�qȬ*? V{��`|`����n��Ԅ��#Qli����@���T�w&ߧ�8ľZ6]&.���߲�SHAv���6��Yb;5Nv~�2|u_H��(|�o���@;��2h^�yY�����O�E�����h�a���n���D@c�>�'@fK;���?�MHP�t�VU�ux4��I�� (�bn�b�4���(�9a�bK����aY�.6��bi��cC�Ut�Z�턺j�TإGw��!�����F� ݤ�n��rs�Q� !2w,F���^K0)NT�BG�G5\A��B�X�ts�������};��S^®)�`���s��^�Ǥ�Ѣ��g�n�x�E=����^�͋�R�&i��IhL-M^Z�:�.��*����v*�2��֙⋝�%�3@w��0��S�Gg�x�	���d�P7yu)E�8\�"��h�`���-�W�Xz�N��H��ZU���-�ĩXõ�[�u���Y6OO59�)3�̺����,{F�0³``f�y��� ;�5p�q��v���fff(�ӧ��M�)G����n�v���{��,h)����j����ee�5h!�'g�a_����އk�*���֋ã�UR�b���t3n��*�����^��2���P�U���yQ3�{IɨW�x%�l:)q	?�D���{zYK;��Q�O�E���,�3]7`��g2=Ø����h̆��h�$E\�[�
�g	����A�S���li�<��_����8Pg�9�SP-O!���,Zъ*S l��#P<>�"����]#���n�h&YE��%���8;X�2$��,�������`o��%=�!G�u�]��fi��4�8�%o�pPQ�mx�n�YT�3���)��8B��[{��,��e�����y����Q���~�5����;��#�ǨL)¸�2q�v��|�ᚑ��0��ڮ��%%�4�E�T.������X�)D&65��M�w�k�9�#�F�ӌ{�aBN��	�����lh�$����oYy�"�X{���޺h*�P]z��Kx�?�:wl�7��[ݺ{��#lG*������q���,�4�B,Ê/�_�E������)I��Z�{��p�lT�����<�Z��(u���Q���x���nNt�C��T[%8,�:�:.���)��ǲ���֣�K��Ɍ�ϸ���j��v��Tm>�;���V�cfu���w������z�@o-�M��Sg{3#�8�V��)ܾ������=CJJ����G̚M
�0йx��Y��o@o:P;M1K�Fa�ـ���ba\	���_i� �c.n<�
�Ƿ�X�����:��<���0��Q���r��!7��>s�������/7���@��I��[^����>O=���#'KpEy�V��|���G
3���`��p�I&��z~�B�l�9�;�Y#���e�8��s��jǐ/Z�*�vU�*2l�f��U�NݚC��G^}�y�N���jAf���f����1ف�੎y't�G���=���^��S��S�[5FР�Z��|e%P^��Tj;K�ᯧ��]%P�+�)'}~&躺d���ry���,�T��z0�.
��o����*�L�v������?Y��E���}@�������ZS��z0P������3���W��*R�8�=|7)�V�ל�pN��u��<�=�{?�p�x�_��q9NLOa=y����;~����2��):�̗2z�c�t��fL,�1sN���?����NC���l��l���U57�z���9a�q/��@wpT;��~� _�Ѧ 8)%ި`fVk~3f��dDzŜk�Q��v�6>������L��j��I֥�� �����r^�H{�����1⅘'Q^�јSe�������d�&o)�&3fφ���N����E�`����K޸�ᵹ`���#�Ie؊�q *��&���ZO������f�>�>2It�=�'a�,�p�ȾGl\�;t���Ug{	 /&f�S�(J\C�)��0����� �?dK5H]}�3��ü�h��O;ݙ���~����Q���a,)Ƽ����)���S����O�ʉ:���2��`��������"�\����
��1~�Rr�Gn����Ĺ����]ٰ3�#��_	��.�˗Ӊ�p�+����<�q%qr2�@7��-g�a�gX1:�t��Mx{�V��캹1KҡJ����r#��d���c��1�n|��Peh��a�5q�a�TOtF}��UAO���[4�8/��AdW�NQ <�Q��	;����ϛ��b_bSx�2;�=��=����c����H�~��H���ơ����ǌh�Ŝ�v[��������$��%'r�|�G������%�������~�����+jqO�n7�k�_��}+�pd�H�ף�G�z	A�Y3^<��>��p�r���յ�e[�I��b�#�I*��HgD���)>_�LX"�S
M;s8�^x*R�읖��Toj�Kb��&�D��R��G&]L��k����nD�70��Z�_i�dG�J4(Im�G��W��.2N�krRxg�� ��3n��h3�)��+9MT}����uFŽ�v�k��G��b�˕�������|`J���]����M�2s&g\F�0}��3kB��Y���Y���lUhc�������6���4d'�9u���N �ZoM[����ae}i�,vc�ل�H�:�Wd��yQ��SM�u�7�e�F:y���j[��~�/���e.���m\-)���wNQ�i$}�6�N]f2`���v��ÞNU�ΥM�|	���rݜ�.���8�{ߺ�����TR���á��c��Jmpxݺ�Aʹ��9�{7��f�SQ<�?H�Y��W�8Ivx��k��}N^Z�r��=����e�^^=#^g0�m����kzz*�Y�5̠{���6��1���nJ�Ё��� � { v��7Ϙ��o�~�	��m�X��Uq|t��4^!6����c�+�|&<I#�O�S�y�x�5��j�Z)�.�Ҁ� 2��-��Þ�(2�K�y׀aCr�=&m��f�b ��lv\�tp�E �`H֪u�Gqj�x-/xk�_s�0��w��L����s��~����#��V����d��1�d�;�D��}.v�z��1��N��Y��q�~Ɋ��{��^[^����>0���|.��uY�F}8���n�)kԗ�'�]��ۘ��!WIDI��i�*�k 1�G��X���3������@���� `3N��횘ޖn.:2�=5N��-��=�u�N&�q=(���w��p�v#�:�t��Ӆ(�8�������$-�l3��A�J�e��J�H����e��/%����+o��.�u<�*ؐ��9f�&g���4*'|�c�U%������0{���"d6�Jw�"մ����.���7/�ǰk	���������p�\�g?%֛+�KЋ���h=͉��R��*�=�:�?R�7#��\�� \U^s��;]sI��.����e�og[6�'�ՙl���9��Þ�5�>'[;�;���:�S|�Q��J��l�vW|�M:F�1���.�r��ۧ��O���V���a��N��I�%�>��S��Hܺ��f�/Pv�x��U5N�J�f�~�?^=��7��*��K�YJ=�٥/��(c���ݳZ��y�E9$�Π���͚�I���A�l2�N^4Z\�઎*�O��
�wf�ݜ&�'�dz�)�,���e�ON6ϤsZ��b����[�NJ�/����ސ5`OH�G{Pc�P�K����1B@�j(��bb��������Ήj�hs+�δ�D��cey\e�^o�0���WT5z����ผpy��y�s�=�J�O�����0��g
����Ř$2�=���@�'�a���i��:�Gp��{�Z''예�ZӔg��+FX_�@�t���dC��P;p�hy���s���-�Ev��j]P��v�y�Ty�:XE��G����d��S�Ąn������g� ��^�3d�)U�?ECL�o5�h��O'����@}�6��o��L�=M�]��ş�_8.�1�QU�`���lt�����k��E7���Fzj��;r֨<�T?>V�qG �������Ġ�7���������I�S����)m��&���˵�(�/o/few<C���Ow`�l �T ��T��wV0s�=��18Ogc0&��:L����s�yvQ��+;�ۃ��&6ݵ�,B�t�1�{��9�9����z���R�--Z�zf���f:��FD�$r���F�/�;N(A��d��ę�����o��OMN�כN������g�/Tۀ���@�W0m���R`|�'���Ib$1�*���~^���~�ݖ�SN{���r��r���'ڶb�d@2�V������o�+l8���j��+
X���Xlw-�I�8��k$�x��# ���8�1���?��Yؽ�1�g!{I]�`��y�_!��,��u�Vǚ�%&X)a�*K�����RB����*��qkOy[�ۗEv������2��� �M��#$�K�9R #���$�fh-F��lxX���q��OF�����6�t?�@�s�G	���B�����Xh2���U����nD�Z�M����L����A%XI��d �J�5/Ϯ�x�j�֞�%����k.�:��)<TAep�R"���C��\wׅ�5I����G����3�����̈\�����NS�Io�3�+yɌq��Gg;�'�.���d�$2�s����w�ҧ�N[��
F��
��6F@bv%�[��Hq�6)�U	�(U��k���/9e��-���T���3%Դf�I�x���qx��6���O��hE��\�I��H$�Q�J-|�e�(c���&0��$�k����q�t��z���'f�g�n2�m91��Y ?�Py7;`�����<�� ��{��b3��}碸�o����nkX358n��K{����*s�,�T&����4����[�p�*����G�/h�Dӎ"�Wu�#zR5b�(�2�w�Cפ�v� �	��t����������G�3���q�[�3�*犬�{�f��������ӕ�6<aKğ�i��s����k�(<�H8F�֘#I~I��`��7�a\�r�k(��6�v�.�P �����*%�Y���s�r�����#l�!�ũ��+4|�\���e�2a��[�^�=$�-l|P.m�)(�&��W�O�;�"�ѩ������vK��i����ٰ��)�Zc�)�F���`�;V�B���$�n}�ВͿ�l���~�'��[�U��{���9���j���ߨ|ÇV�Y���.�5�e�bމx�\Zf�{�I�'��sG���_��ư�p(��v�G�y?�k�t�2Յ.7q�,v�:ǿ3�x�`|l�tbF�¾i�%)!�y��(Sq�b"���{���q��35K~t�d�\��K�8AY&������E����:1�E��>�"O��Lt5S�7wd^"��kƙKd�����8�U��,���ާ���As����sz�Ň������� @L�sxIol�8������ 1�f^i�Q�T�m�Q�����y��=`�H�b���ߺl����8���"3ҹQI��j�ͨ��}�2Mg w7>ts��8T�����:�|�	E��	v�ƙ!���_�վK	�i	vfn�qO��6�ϰ"����6�a���F���;=��ۀ$Y5��H&�e6�,�@�R��@��gjj>0��׌�"c�&1�F����>���DA�ؙY��Wpg&n��:���NR6�7�{'t��;}�"���@���JQ��܏`n/l���&@��[|U�D�'��i'�{��\R��P;���4p�h�Zn�ڔ:�xYŵ ;��f����uLw�?�j7ʋk�����%����P�WW+�	�^cX�*��&�;��y�&�l�YA�O�q��[��A;Wv|E��f��m]�J;�ҘN�Qh� �r�<l���X0��q��X8�Ý�"���êbø���|����"د9��^DbV��%0"�����30(��nY36�L�j�;�s&���hϪ��6�	v��[7��7ʽ��9K���Q����.�p��0[ƧNzС�Gu݆�L�7��m��7�Ƥ�Kǅ�I<j���R���{��m�q��+�}�ٷnz�> 7�S��"�i f��>Zw�;�>��W6�sB؋B���S���	�'0���%x]���{^;���BB�%�wd����
�1g�Ʋ�6��xG<�nc��:�P�M�`�,1D}�1K2�l�T6�p��� ;�����.�L�� �i��iv��v���?ٺ{��v�4N7���p��@��v�؍�}�����O��ôF��L����$�۸��"�6�鰱@/�SD�l����6Au�b1�j���Ǻm`�7��`J�=v|����g�c�����~��Pۮ�ڎ�"�3�39�ٱ��������wo��(�����:g;A��*�8�����2.�.��l�dl��n&2��6��q���0 �A���;`�c�z�+X���&���`*�b�G��i�`�}��g���k��`�N<U;�gJ\7�>���	�o��ؙ���IJ��q>��0ݽ]�����̋��F�'�����t�R��qb�EZ�%1�ץ����Ɯ��R3�cp���[��b,I�!enN�Jv���QU{@
ՖV��g���"�g���yFw:U���g���8S�`F�>3�{Q7�<�9ї����k�.���n� n�!1.��G�6����n�2v��5i�
tO1�EQ�R��=����g�m��&@}��2��?J���׀%$�	G�)���޶����i���Ơ��i��d�_k��Fh�{ԛn�!3R��2�]<���z�8f<C�ٗ�x��/s���`�͠;��0^л�d����4�=��"O�{<�����K�*ٱ���V*8�����`�x��G��]`ǖ��Șiۊ�	^
&[��jۅ��Lj����q�E>2��^�Q)B�^q��(fP��L�����e��������q�glw99�9��LGPi�<-e�+��6�¬�(��6�'Ay��lM��qZ�ˊ��2u1��oO�\�xm�=	�o���3\AX ��n_rC3T�v�1M���b�ԵL��I���%��q��{#B�	�� ?��N'�Bv݊�������-@�v$��D�V��N�>��t��0�Fs7�6a&.8'��ƕ�bo����Ы%y�b�bG�= �}��.�|E�����7��*���]�	I�SZ����Ku���Y��碞Y���tG�7= �KF��֍�ǳ���W�%�=�v�x� aw�9�]c�JRLH����i�&AZ�R�ļ�ƃ6{�bk"�)�WY�ͧlX�%1i�.�^«)5��,[{z.]�~9t������#`W4���j��ecήj��GV�۽{�����8͊D[�5|U�G&���>��Ǟ%L蹸�p�{��Q��GB�P� ZP���Y�GE�-��_�0��#���� (������l�T�6|qP�� �����g��7~W����#�nĐv�w���ׯk�9��̤3��Hw�}�s���ł�.=8�b���/�yw���u~}��˅�i�<s���14]�h��J�j�T��NQ�[�����l������]�|S��$Fv��%����`S�b,��Cע{�?����1����6�E.�T��2u5�9ӎ��������hn���"ļ�Aϯ}��Q���e�GM�{Ouw��Ĵ�CAE8Bm�X'2�&�M�g��a�27��P���l�o|S�z�͒T��LbX�5c��2^���R����]b���Y��8��Ul3�JY�*k]�V��O��}A��/.��"lQ�k%�H \�&؃<�n)�gD5���0F9���n^`�v��B^�[��G����H�Rc� Ř����0�|�"m4o^*�FL��DB�0��d�}�����8�VZ�H��U�6�J��kv���c���f{E��*��y 8B�F�G�&�]��t�uya�Ȑ3ۙ�`;L����̔�`%_�T `ˉ�!5nO8�q�8��u��ԃ������M��3��R�� ��jT�\�=���;V+ut�+����ا�aǑ�Q��#x����DA]�U��Ff<Np��l�3d
�/Cu��t��
�!c�8S��nx�/b�H��)�gF�a�Ԡ�u�Kj�y�rP&M"���0��Hw)�����<Ss�G�,�Eq������p�mU-.S3y�L�]�R��wd����}Eu|g�F4o�@}�$��~�L,gz"<�:W���Of�#�(�LM�.���)�-�Յ?K����={�QD ۹�+�'�b0\T\g�Q�������ͷ���(1��E �8Vic�V�E�$�����8��w�dk��Y�|.g�KMe.oF�Ϡ�Ay�ƃڤ'����O�n��f?d$��8���6�g��bs��,��Ȟ���;����P��l�Xq���kQ��|��?*�3�%\�3^\�����Cbw�E=�^S[�:��͒Ju����<%����ư|��
_Q��e��~3<���F���B���<N�2�)��H};�6�N_�>u���6��+�<�hJnpyw{�	3{C��~Km2���a!(�?���G���0�=pý�F {��#}�5���)&v��ij�>y��4~:���jbD��m��>����>�[r��W�S�Ylwq��[z9�~\w�u��k .D���/��X
�F�W�d�㶜<7���a�g�϶[���%�2�2�f�~~��W���ōh�|O��ڵo-<l���g�";B!���x�Uՙꮣt�Y�p�:��S�;_&�6w#����	3ۙ£�ރ%2�^�)�NL�8�����cpkX���:�lS��C5�I��c����=u��v�$ �Ƣ/����n���V%?�"������V\[s`���!�gܱ�<�>��Ё�Z,���δ�;nՓ�,��h���V,h�9�iEA�����x����d;�2.�z���a��n?6�sm�=aKr�=��/6�M�D5��b*�9�ׯb�:�M��n����M�Y�T�O�~u�����
��b�o�q�Y�K\gߺ�	{[d�p
mX�������}'͡������
�Kl�J���F�͗(7��lwuSB������{�!�,(T�k#��`{�j��¸e	n���:��4I���ώ�Sa� �����2p����#��(��f�:�E
�|Q��I&�����Y�O�:����t���3�iɁ]�!����W}1�5E$;x|?��0N�VU,K�il�j��e*ZB�i�
乲�p'�1��_�|��R��hɰ�2�7!�K$�3;3��36֝�悝�t�1�a
�m6[��:�����JG�Wc�L#{�9 ���Cm�8L\��T �[Q�o�>QG����K6R0�2�rX�����t���o�KWG58Xw���:����k>*L7BT�⻬�E}_�r����߼��ºh�D��x.����-����̾��$u�)��zc�ǝ]o�f�׆-Hu쐙��FQ%3�_�v�$����I;~Q�T�Dhg�^��|��c��'�O�ΜhXR��d�yxݨ�`Ok\�Ӳ�G�D��KrV~����V/�D3);`[��n�����
�c4 `�,��?���]�*�^�x�]_$���λ����`8s&�V��1�'���x�"�g��x�Z�d���N*���P��ǵ�*n��ƒͿ���S�n\O2:�S\n��jT�0�����O�b����+�?=6F9VpY��p ��Y�u�#��N��r*:-����x��D��{?�G����ǪBO�2s|�Sw��0Ml4�1�f��SgzF����g��=�����<~&�)�g�)�!+�WJ%�Pm��
Lm,��Q#r�7�	�j�4�.sVv�fE�2c���ؘ}Y�]+��<���/*���9J{�p���f���#��~t������KwW\<����[Yy�`r��w&�_>5��B�Bk¦��&e�el�<6�ǳ��;U}��ޘ�ƌ�?�u1L�Q�
�����q�����F��ߜ�su�}�{-��T�Q�	�e]�e+=4��X�]P����ؚ5cG�G|E^Wse��l@~̙f�����Z�"�Y*�3��x�7^��|��p2<s>�O�f��cOy
3z�]e���
auQ��c���zh������b2b�l���򓲀�0��X�调��W��TFkdd��'4k;v��c��
F|Y�9���M�	ux�OT{�nV^e���WF��U??
'�����O=U�G(��G�nN�1~Wd81<J�CڳT���l1S�f�=��"Cf���H�&a�]�I��S����x�	�=�)m��N�#�l�OZ�:g9?]��I�0��3�v�.X=R�k�q����Yl'	�Gn����Ǒ�%_���F�/�'�� �?{���1�0'�-Y��k��0��B6�j�����X-ߍ7�`H�ޮA����P�����iZ^~��O}�
#p��SO����ٰ�e<�'�&RJxr���K>�,I_��ݻwcsي�����w�`7w�g����"��F+���R��Aڿ&�}�;o���`-ŀ�1O8桭��w��ˠx)�΂-��@x}�QF����RIiRs���_
�
��[������#1t�}������*x��P���	�[�VsuM�����֌!�O�( �S��9�b�,��̚���D;���c%*�}��p�~����*��r��vt̒�(������B0��>d��:���<�Ý�OVY�D
���h�\�C��V�q���p3�}މ�4o&�L��{qO�\�M��rc�Q�/��f��Ygv���/b(����� ��<���@��L����h:���`2�j8��ԅ���l�����r�Cy �]����m��gö^��)1EI��F�x�����P��	7G����[���c��o�z�y��m4a_Ѭ����kz]M���n_0�{ �`52u%�m��l�4��	�g�т��/�C`�G��'���;�/�mfim�q�=��t����f�X�`��M�1,qdM`�QkQ���<&źnǙb��P�6�n��%@��'1�ߜ��;npf����b�8�p�E�d;�L��`d���3gf��Y�?�Rc֙�fC�'�l�f�+�O�y�{�T����蹯��@88?<.k`�����ݺ����N��I�� �h�oسn���H���v�<��W+����@����~��޶S�t�1�w����9�q	�>.Ѥw�e��I2D��0��pô�Vԫ����N���C��Lw�)�4�j�r&2�l�wn� m@w�7�H��P�Sw�����Xh9�.0S���A��ƹ��>HN�P͛{���R2����(��.��Cuw���
#px!��,��Cv8W�/.�*gL|�lZK���U���ʂ��Ә i��	�/�mNW�H�n�z��y��p���*+���^
���p^���ʹ���o�et��y,�ڎ�h�^��=������C�<�K�5`d��>nEu����S�'YQ̭w,���~�p,w�xl������ں��՚�����r�0���l���`M�Ϝ�D"��i���Y���nFs��/{��o��ܛ�����@p��[�?ww��}B�uU�e��	�-}�͝���G /�y��d@�d6dM�*�p��2�PTE
��k���P/#���?�'�r��v��o��]�8�@B��U��U�He�&3`��5���]��)���Y���N�}�n��|��Dg,���W{_�[�U����J�`�S���?5#a}nf�&�ɂ�Ř�0IGy���������s�]V�|��M��:h�	=㍍�*s`�?�~C������".*�����½TÔq��W���>�����_~jp�(��(���_>��R!q��T�T�V���ͅ� ����g�}����NS�X����P��-�p�Ν]�4}��^M�U%�����%f;k��@o��w�܊��_�N]�� :�����N��[z�����Uŵ�^uPV����ȭSp�R�v��Ա��T@9 _��Țݭ`ȃ%duQAyQ,�'�C��a/�J�y��Z��1����Q[ۗᆻ������)�~�t��}A�<�:�:���8 )fa'�O�eY���(�
3/�Ӵ�@���&��`��[���4�~q���j�[-��\(0.��Z��������G�Z���EY�>G��'j!i}���k�����)�� �}�ھ� VF{ln�����[�R�NA�=u�g3�1����c��%f�P`��ST�!K�n'�K ^B1�z��-��2�{��?/9ڇ��C�l�\��4�e�z�cI	H����F��y��� Bbs$���),��:�x"�Pw�9?�!���!�k90��;�`�lp3���pA;򼮎<RK��(3��*!����%]Ӆ�kV�`@��� �8�a��,���BЙ���F��|Ò��j�Qh��C�"�_Բa׾|Ɋ�"�4bf��/_ɴ�tk����v<b�2�Ì�vV���wUm7��Eg��S�^�,}ŻPZ�Ν��c�[S�b�(�4�u�&���yd$��_��Qb/Ea�#�!�c{�o����~E�o]��!Kp���|W1:�!,�=5��%�YM|\�hN�'�0l�T����i���~@� �X���*���蜅�e�����DZUAڃy���cd�਀�޹�f�#�c��)�n�TB������R@Q�|�����6$f7Td:�^�SAE�w,�'���`w�m<��A��W �yl$0FhZ֍eEĴ�c�4���4!$�7H5�p~�n���5kǑe��\�+`�OD��s�F�X'p-��psl��������D�=u/.}��Qb��b�������H��)]���ZU3k��AЋ�����E�j�s���C�Mv$�vaD2�=�X��n�9H������ G�����Kۨ���<�|{�`;�kv��d��|��>ހJ�@�-�`�.���~�8�|;B���s�<���#��R*�����_����HQ�Է��Z������P��dҿ��t!�o/�*�y,P%BCڠ�^�#˲��ïI��υp��*+6���pT2�Y�����ֱ�5_�?�f�?k��M����q�
|}}��	��_V��6{6F�= -���>La$Ōu6��6N�-� ��R�'{ �gI$?ٯ���R�]�zkw��`|�f�����x����_!����ƹ����!mxΠ��V�dG�q\8֒@���x�~y���3!�$
�W:x_Q{��;���`��8�<�f�^��ȑM���W�c���	���6X�uoTsrDg��#�%d��R�Pr;����|��Ww��(���~Վ�����_��0L���Py������o���Q�*����T��_��>�_?��|��U���!`��:ϴ$��k��vd�X�nf]r�9��w�������LH�����ܦ޲~4[�<U�d�:���#�K�)ƾ�x��jsZ@�C���r���[Q������7��s��Q�+=ZPb�������pw�3���G�������a�$��r�<�i��td�,F��x��5di�]Nص���M�8H}_1< s	_M�Ȋ:u��"���B�Z"�w���^���d�V���o���bs}�uv����ԩ��iZg�/�6Ru5�3�W���D��������!�ȇ�\����//?\�4gu>���A���Zq�����M+^�3ý�(n���Ac���a���.�8r^*�T�}�N�H�aT�=U��s-(̪�w���:]k��x�SK6�?� �g��q{( �wL�)h��7����t�tfH�^C<]�g�˷SG���D^^¿�o@~��M����|6/���޲���8�Is)H�@nJ�)z�.'�p�ۇ�~��ds�ݎ�h�WT �V-|x��3�	w �7?����Ά�%�D����%����y�j��L�u��,%řNBC�p�`����h���vdA��]�n�?�.�,ȎO�����T��:���������R�8�}]���W������G�ol؉}hHv�	����Ə�}A���J_�����я����(C=��o�� �yg���Z�1�(�8�_Y�TD�7G�h�Qx�O�ĄEҡo�e�"����vI�_�{���f�QPϴ�q�ڞ����7>p��������?�� �Ah���t���!Uk����*{*3if�{1�~�(�xo�����	���[B�@�b]�#h��v�׊�p(����#�8��H���̈�PF\��N���H�-.����=J�_s]g=�psۡ����l8��@��ð;hV�t�K�L�4�<<Pf�����c���6NI��F�C�p��Cb?*G�n�H���m���m�g�H���� �p:�xAG�?�S~��W��.|`�jV��|0�ݞQ`�S���/q?�ٷ�1�~�Q�{���K��)I4Eq/b�HMk��!�L޸e�qI��?V�} �y�ŵō���^{���[?��Pǌ�����;w~t��[���;�5<X;���*I�s�]�IB��3i�"�����.�gd�K3'I]6�����7�:�a���wT�!lz����ڶ�n��w��b�/���yn�-'���v�᪗���%C�R"pY�KC�/���}٧�P�s
9/V4b���y��jtP�K7/ʽLؙ�!׫�L�e����R	�.)��@�u
��[g�>���x�����~����nyܑ��1�SsZ����mEm���i��P���O1���ȞB��RQ|��)��������^�#��^$�-2�cP��a�|/0ogoqL$:�:~�ܪ]���<C���nR���[�����ѡ��7o���uI�Yqrg^�Lv�%b��aM�ظh��le'*�E����`������[l/��37��`/`��_���J���~�
�����5�o�Ɏ������?/>�о�������S�� ������)��B��PG����裦h���$�C�u9\_��*���/���
4:�\�{M��V���$�� �7FX^��gw���s���ݻ�j$;�!�����b�ߞ�
��ֆ�@6O"+�-@�9U)E��:���\ڑ��fO1�39}�W�	�K��Na�L�#�g�.)4<����Vר�F�h'[@J���'����曷�y��q5����{���׼��w���tt$@hBR@±Z��R�G"�%�'ٱD��\U�QʊΙ���޻E5PU�'́�9�Fs�y(
�~0Q�m��Q���#�� N���O�K�)�~�m����g�V�_E�>�thߖ-7�ZUst����r���h��f��p��-���>��(�tV��"
p/����V	[���¹�~N��� �QW簸gP�1ky��������B������~}Uj�5�0�Ic�}q[�/����hyMM��?t���i;�Wh�Vl!V�\�W3َ�bC&<�no�bA�����_�Q�]"�cX��]1�lY���3#y�Հ=T�z���630��'?�C1Ga����뫒� � �'v2�����w�ly������f�<P��JU4U�Q/R��u2���z��v����]�[���?���ܺ**m!i��Gv �%%z	--+  �\�h/�=!�K3[Z��O���+�7���3�R��"�;w��|��#��C[�ly��������r.V�]�������>U�
�_5Jb"�fh��$���n��Q���q��?��'-�i�׫:�<��JR���ֲ��
/B̕���W[�����7v1YЉ�]����<���W��C��~�o�;Z\s��}�R��
fv8YQz%�����Z)Ig��$�:��b�w�Z�ǎ�x�(��4,�'��j�;�^it�䖒�䅈�/�o�G���ōP�7o;G��W1��#�;��+?Bg�|Շ��<�&�My����w0��@�� ���"VzRiN����v�]RS:��~ &2��_���գEC�]�#U�>r:��,�T�f��N�� �zq#1lE�sӑȾ��}�<�}�JR�f�ok�������T�1oG�Q��p/%��E���
����0��@v
ꢦ����Ǩ��x�u���t,���dYx���9SS��X���S  �h�����a̜��8��'�<Zq�3�r�a��p����V�ܹ���9&3�=S���A�E,�t����6G�!�!�DJD�E%�`�0�f����5Z�(�TWQ�xt����x5���NG��(���e�|#|�H��j��m,.���t�߆���7]�����v }%¾��m�W�n˖_����C�{�巁P�M!�̪��OEm�PH��Dw�E#��dRM�[-��iuU�M!e�:�Q�#J����� �ʚ����Ӏ;g:�AS�,ug7��|���)�7�/�}�J�vxu���G�������|��ܑ����]��đ��є_��+f�ң2r�ʲ�甬��"�x��Da�=M�)tS���;6���Q<<d�� �jc:;f�a��9:�����3�>�,���%D�_��/؟���c��QdnX�ѡg�۲�w���)?��jY��\��Ϗk	��L��W�t@n��j%�d���j6{���/X�D޺�?��Be�*��wX�qG$14��!Kr{^(�ŗ�.�X�������3�Z��B�n��a�	�R�N�g�w���o8T2����_o�Yu��gm��� a�j'����X�Q����������e�!���[K�-��N���H��M1";
���Ն��!JB�#y���p�?}�9p�c������f�~��G��
�Z��y@w&�D�C���ξw�����a�p��Z���;B�#�ET$��Ea��R)~I5k�����/��:��6�>Z�e1�u|)ڰ&�Σ/�K ��Rҹ��.\w�矏��g�����3���@���`;����|��?_��;Gk�|��Ý/��dGB
�ٍ8���,�-�����1v�?�b�=�����{�}��k�%����F�E�*.V9�`��lga����z�>��+U������z������~u�>�>E��;��P�s[��n��?/^�s���i��NR4��	%�'ዟ0���W�}��`�b|���ڋ?�?����������>|x�ŏ���*m,}���͐u�t|�������v&2�1۝��b��}�*�χ}w�|]���8��J���쒔	�0�M7"�Á;�, � ���@ɾ��$� >s?�|u�5��bm,���
��k��-G�:�d�\Ͱϛ�G*�V����C���Ζ7(&���gÈp`\
 ����EV4�Z���x����Pp�s<���07Ȯ�
�s���o�0'�>>����~�UX�d�~���l?kf;⾓������_myd�P��]o�2GW�j(�q�����I:M��_��3Ȋ..An~���3�����S	ӿ�����T@���q �45i�ʫ�n��/��g*CJCF��-[�=�l��b�ղ��I���9��+�َGb�3��F� }@E�ׄ"�jVMU��!x�)���g�66�����*�_܄�a�J]d{���.�Hv2e�Π-�)�-��<������Tɲ��(
�Ҡ&T���=���:���q�tG���q��7�4��BJi�2�I��aw$�����2#�g���#�~,�/q�r��=V$1���+o �њ�E9���|^�&��/\�s�{.�s��Q������@�W�xN��*����ڂ7@���H�8�����~�+��Ɍ�����g�U
;��J�;S`����3|oz��_�UU��&R�x��H�##�D�$.|��v��J�����>�����$��4��Ѡ��
�3~�j׵��7�k�Ȏ|_Ɏԫ���&��{��ev���{��w��{��fqy�;?�E��j����j�Вr�:G@��'g�D"T�I5�� /���6��*9i\�w��q��/n���m\�W�s*"K+W^�l��M��s�븃���оw޹�|��g}g��{ ����&#F��P��ۙ�'����'r�%~R�ك ���=��#ꁀ����q���|���z������r����N2���G7�v�͚_��T�恞w~; ��IV3�P�@�'�v�~"�gf�Q�7�����TE�Pl��� �5)4>��ޭ�6���	'��v��*��v��v_���7���P��7���`�����}�kY�f7jS^}h��XK��v�L��Q�(Sa\`��c�3�1l1j$^�����dF���.�ƔӋ���n��6�*%H��4�B��D�(ƌ�^)��Ȟs�e'��mQٲ�ҏ�s���s�=��t ���)��d7���9�qa�G"����3�|�Isrm~���o`9��(	���)<Bv����	������>��2^�beg�>nR�2�������An(f�Dۡ_�i�֘�Z����w/�;.���:� 0�!Vg�D]"Y�a��e(�:�l��/sC�{Ԓ/��� ��Y�mV��m��0��:)��4�<C�\p��S�2��/^���y�N�?��݋�"�E�I�>����̇'I�s��f��6�'����e�&�$=5�n��A�����Ef3�Z.���q�cʏ���J6A��W#^%F�T�����.n�^����8��24��x���ƍ7�8�)nZsx����SP��}���R4��n�k�Zڲ[�����yٷ���ד���f�t��qР����������[n!��.�C��6�M���3}��y`�W$!M���a�e��ke G��z���(x2�x+�������{���r�f�x�(3�&'>��כ���$n�2r��q��K��cHJ���'��I���p�v�܀�����P]��
LM#Ҏ��u�{�ɟG��;�AG]��4��Z6"3�D*����5¥\���8N�ܝ|?�[C�Z�ܧ���|�����ۺۈ�����Jl��5��}��!�u���q�8OK��\��#�
C�cҫh���B�j(h4 ��&pe�؜�V,��D�x�M�i�@-�o] �D�y3P2��lm�K��pE��&۱��HP�C���''݆�i��`���S�
F����4���u2J�2�b�&s*"���*p�]��M�jJ����m��[�P��{���w�fR��d'��-���D�����M��oޞ�0Í1DFs�t�����L(�T	�q�U;P=l	�gql'�i62!R�G�f��T�ŬN4ڕ��I�������E�[�{T�|D�=r�D�wCYP��1����;�"���ɵC�᝿IK���s�vŝW#!��g�lz<���]/�Q�ѓy��Qm�9�|��x���O��42Vy�J���t';�?^�����oyE���y���SL�Y��%A8a5�;I�gq7�Doˌ���M�ߘ�}�D�6�j_v�����I���N(����W#���F$X�R!���n��*JC��r��g��}�b�������s�eJ���x[l7��T���y��]��ƀz�c,
���0[� �����5�T�����A#���q���Yeb���5��LD�W�x��>��R�����b����x�7htT�;V͸��%PB��������nPb���;��\pZ������#��[z��ol�>1[ ��6j��o�X�û����w"�bH;Q�yP�:��~{p�xz�]�w�� ��8�V3������5m���U�$;psb�wM��q~�DT	�/��x��<�Ŗ� �'��H@>Ab_������+d���n=�p��谖@��x�BC���g�����JU��1ڰ皞A����-�A�w �T�eL��|M.�Î�k5���4��!�&svO_<Ŭ�%�����L�� �D��﫧�v���Sx����e�������X�_��+H��������x�{��O���#
�˯>�s0!�b�}��˲���tU�e�F�]�P*�+�������%�'qr���0�7�Y��F+�{7C��	:귷�Q��������� 7���?�>��_���xűi"��6\������w{�pf��Y���f/�ۿ{ɞ�)G��R�ۂ��Y䳙�����op$ᛘ؟n=���IG,)C�On�J�ܼi��d<]5�,�Z���u�}��-`��?<y�dwwwސ3�w6�n��x��c�F&�~��Qe�KM ��a��8�if��>U�kl��M܆N:]�8�>�1u�v����-��1u��B|r(�>�/�C�M}��T���S���խWo����?���>��헻�S�+�V1z,φ��Ü^��ތOjpU�U�?�]�9��:���	;���W��+�����gG�۶P9:z�x��n�����!�9��\�1�߇�B7T|���-@����ӧ����u����x�eo��%���:S���q��Fl�������$)�e�1Lz~��3���T�"���^�܊��H@=������������]æv�=�z��������x���j����"��è���^w�nG5�ztӪ$q�����/�52�{���Ā��؍�w�aC�P5ʅ��\� ?�(����g0�ހ�[��[��>UF�>x��a�[p��_]�u�֭��Ǐ�������!�۱��\1}�׮9������Fcda�a���N��S�p������w:U��FvBۼrE�O�Sֳ����� 	��u��o�4?�x��C#����	��v��{t�
]�ﰮ���/�`�����9�ޥ�S�="H�������ks�?�,�~�;���7;�?�'H�΅��<����T��Ԕ��k@�5�z�X��ǻ�����pA{��\Go�r��� n�ӟN��������g�C�-�E-��b����{��0��	���>Z�+v2����w. <
N�hn@>�b�X!�>���ߝ����$��ߓ7�oк5e���g�$�Ϧ�	:D�:�;���uܯ�����_~i���?�X_q�:¸����w\@�;\��]uB�����.f�{�:�v{��״���ndR�L��q��������?]Y������7:��:��8�*��l���y�j����c7�V&�,ܟ|9��?��$;˲4��:���T�����{/&���~TaGm����� �|��?�ۛ�W@ ex��,�M
 �5lsvS�N��9�7�l�\99�?�/T�����pP_)��	�v8(�i~��ǗO@��*�V6 {�fKj�M�5E�@�:�>� �]h�0�nz�|�U��cB&����9��NO�5%����L�u�x��{}��o�Zm�&s���lVg�c��,U��p��fd����ƻ�v�+�A�v�frM>�m��%'M�!���ygv�m�e�9�Π��������3͚+�(�-ՉO6�:ߥ �����
F�������+�Q� ���޵p�����2�-Z^�Kb���vc��(�J�rJ��<.>Bo�� �V#�w�ߥ�� ֖
�}�a/x<;���;��	 ���51>D��V 2ߍr{�A,&�a|%��o���˦�-�fy�ؔ<�Φ>7�:��[.�U��N\���ZdG�jC�V��ņ�QY6@׃M�_RU����P^�x��Gl��:���}.��L�-�<��8�S�f�Vk6��K�i�1ҫ/p"�cQ���F/fB���݋4Z��XKn��-�F-����!�h��DQ��o�[ꋾZZRc���2堚�N�k�%O��	��k�"���j���w�\f;�Ԫsz�a�D� 3���w���zg�����d�a��֊ǍNQ�P2o-�}��2��`4�(4��?�a�ICh
�����<�`�6����"-�� >B�Xܞ��z�.�@�D��8�V��e�5�	!2�勑:Σ6�X�brco�t  g��0��6B���X�������AGv:%��!�#g��Vu���'�'���ڎ�/k ����cT�`%܄G��� k-�]���.z�e��͢�e�����ƀc�e-T̺��D�V���b��L1��.>�g3xl�!H�}�����Bx� �ƦWG��ӡ�� ��=��s�{�f���"���eyL�Z(Q�L.H�l��{`�ΐȅr�L7�� �)"`���,�),�"�p��%��(-����T$XLx<pl)���2C:�����%j^i�Eu�'m��*moi��k�Lǁ���|�N�*�3�����\�	�����c;c5��FM���t5���K���^�����-�0��+��N�T>�_� D&O+
*�����Z-���*{�}YSs�Z'-6=UU�F# �8�YY���a{hu5��4����a� �&�RS���X��tll0��vv� �'�0�����1�50���T�F"N� Т����q�4��-���ۈd�Ε�>���y�R�Yp�C��7�:�z8i��'�f�ŠfB��g���iQj�L��{��?|S��U�@h����9|iŞ��F}�^���|��O��S����oG��I�Lf	z���Ug]Q�R&M)fkW�#����d{��e�98p��.C�@ԓ�ƂK�PY�$YQ'N�"�C;u:�й�`R2<���S$�>{�k$j�Z���i!h5'����Ҵ��7MN 7xp�A�:*x�#��իq`��r�
�N�Q! 5��K���������vw5��q���.�rT�ீ�h�\�	L����8�jHuL\��"��8���%#���7����N!�) X��p&�)�UP%��}�+�����͐^�Ǖ��!M�ѐ2Uh����d|�E�/��$〛��AZ���nh��ɓ-:��<.�� �و[lO�sٚƶ�rA��:�o@|
`�,�ͧԱ�)�{�O��%�5$%�J��7:N�#-n�+�� �G9 v�X:��;%6���eh�� �ʡ9�� v0�0F����?+2����X�
��>z��*FЃ��+�F��u5�,�	��z�Tu�$<	�VU���V+	/���̈́�d{K_�ժ��-5P���:��Y�� !H�`Ďg�"S�4�� �o���q'�.$�Ž���F��#�yR�X��&�޸�O]as�l��F.��ō5����fHr��sPuE���i�	���H`CA]o!��m�L�u�<��"�%��t�X#z3T� ;,$7��Pd@#KE2���sX���d�0�uk�XA�_��f����?��Y�N�6V��/#����@�s!UK��M {`g|C���k����u��X`9&PG��#"�y �T��Hx�N�u���,'8��פȴ�m���������2���YO&��L_���/���@��WGv�v��^��X�h�\�}O���if��F�J=St�T�Zl2�<�^��Z�"���@�q-t ��H�V=�l#�YȂ	d����Fn��vo=�����n�g��D�<݊��5�ִ��e�;FG��_|{�ܢ-z�o)Bݙl�WW	$�*�:8���Nv?Q�
P]k��1Y:�AP�*��:�4�X�h�Zi�S�jh�#� |1S�����A=T�	��.����:��kH}>��{�y��C�G��<�W�MM�o���\,֪�<9U{m��[�x�	��y��l�qet{�^�k�t'����>`;��B�n�V�<��]�"��[�[�s0�A>�A��T�eE�@_*&j��jo/�?7=�y���<�?n���48Y�R��Z����[e�bUf� }�;��F�(����jd�NZwD��#�R#�h`Pt.2�V���b��q�pD�[í��T�\�j��K佡�6Tp�ebc��&	Cdo���Um�C`�3w񉞋�9��G�/���ݺX� ���.@v�0�cIm5���\�Kdyv�x��߾j�����<H��������-��=\�S'5��T��R8L���0��G�?#��9kKe��e�^>:�k��Y~(�� �����Sө���~̮l �.W�ug݄��:�.N�f3���:���bhv�
C�)�/�-���@��J�&���.���t�,��W�{���T#`�+���R"�?�A�M�A��f0M�7#�:����*����Y�l�E�P`%~��3S��2\�����!�w.mg�5�d���Ů.�v��g��VuA��/?}���F�~��^sw��7�֋���~�D�h=��rd!h>�6=h{�az�Z�eBNEQ����7B���֨�?��V �gˑ�ǹ�ªKh�3����B��A�4mu��2�::��~Qd�GSb�S�[n���Z־��)uzV�淥�ӆ�<V���Y6`� �l�l����P/3b�|����ugP����'rH������4�^%�"��v����o�!��	$�G��Ѳ��O���o�<�bh��A�R�6��շ
x���s���*dzK+��a�vv��=�����vlīClҘ��;j^ۓ#��n�1Q����2��.x�^�1k�� u�����H�A��+Z슗���	��2z�%�S4u�1L�~Ɍ�R 6��l��5h�����[�']M	ٱZ|r:E�`-,���DV�ө|J�ڭ�nG�+����<�(��-Y饴̨���u,���I���lx�&ב�nRv�% X��Q��=�0Q+���b���3y>�W�Nuз�k"���n0����4��R��=���M/�wK�w�!�L�*>�|�w�NV��n�n��gm��a���*aY���W�����M�&�>�/�W�hӥ0��΂�Qf���^�R)��#N�4&E���+1NUe��n�=p˱�l��24cc�XA�h��r8,��RTi$�۞'�6ăRp.���@{��LIJ�(0FeS�9��#���h&.DJ����1���p�L�	�Sn��-��� �)3�������lÔ�ћ�H��+�2�P�6�����X� 
p8<�Ф^ڂU�w|  =
S����K���xF:�	���ݭ��F��簛�cw���)@O�v�d���9:��mV��c��մX�K%�9��;o+x2�5dN���Ru"�t�&wd�r8@��_G}6�e��e|)G�E���
M�0*t5��C����T�`��N����F��?��W��,�H�-t� n�((����u��(t�9�t��Q[ލ��)[)'U�%ˎ0\gJ�Ԡ�e$���5��/�;��N͖8N<�_?�_�S�.���e�����p	[��ԕԬ��'��_���v/�a��^�֠JXt����~��![n���l�����G^��SFtA Jr�s���ՎHQiE�l1b�DM<�0Ur8
LkL�ڬ�*�@�N��%�K)du��(x�퉳����ڱ(V�e,%nF9)P�w��ЂZ�$P�J�*]!J#��s�������$�=z	w�CQ�X�ڙ�?�8
8J���ݠ��ȹ���'RZv �@L�X[j+q�������8��wPLx<�4���\�ӝX�K�P���-\�z��Qogl����jQ\&\Р2%s���f+��d�.皇��vΉ�����Q����t��;��?���\f;V8��ȝt;���}�|�D�q�?�@���^�#qbZ�B	+A|J�؛�o�5�I�t� Lv�*ۜ9��[����*S��h7m��������`�;;�N!l+�@��i��[<�Ŏb�$2� f	lU����g��� o�EՀ�te̠i��~����
�`�����~�����<���ʌ��N-|��/I�pY���r	Z']���=��ihF>��3(�,}���{�=m��R�ٰ���/�=�тح�a���a�����7�bg���v��bv�L�'&�{�n��l�[��S�{/ȌI��������EF��v�����v�䂍��*SǇG�6�uҕ*W(P�2�x�S�D*��� 1�iTqE�f�N�����c]{�a7�h�?��ڱ��x��.��+������Z{��W*�^���v�:�W�*�n�ݞ����P�!'����	�]��;n;W��ҝ������'�uJ�Y�'��Ub�����*Qa��T��&�]���ފU���.��c�׋�*��q��c��?>:j�p�n��Ad��ȇ��g�v޼�З�LbW��A���&bmh٣�B�V17?O�y�I`��#�{l̑m�/��Ug����tg�tP�O��WD��G �h��s��Ȁa���F������(J���<t9�:�u�G`�\���7~�毜�- �maO�s�J/T��۱qh��*�s) �5�t<qd���)�a��&���FG�{�^b���չw�.2[�*�����w������Ia�[
B!���������@X���i��ȝN��������*H8>`;g�e�&����
��`��q"�qc���a?6~V��	���I��;�����ӝ��X���0�����	��c�����ŅY��搚�~;�_A~磏���~5�O*t�����̛ŃA7�:�Y���S0���������Ӵ_<��m5�(p"��8�wF!0b�$��,�����g���gb",8��FWv��G�	p^�)LI��c%�s�����^8��������ly�|o�qO~������+"�s���I.���,��
���ʼHm���,S@m�<�@���j��a���џ��p�.��e[�#I�33���Cp ip~8I{3��!��a\��hU.����7{�c�µ�p9��5���Ž���⛃���TE��)��0���s�|<���V��n�!;�+]�[fˌ�򏏽�{3~��;��5liL:5�q�e���^
)ZRS��iJj��1@]�Ͱ����L��9�8�W��jx���n�VPY�t�oV��(n��Ąo���D���~��9J2��-��\of�?�v4�l~j�ρ,i�ٮ'	�6����F�?Ͻ0���e�ʈ���%p]*b�]sd)� �_��e�	G2,̀��K�A�e�rʈYp�fH��*4����\��(6֙ᨓgGx)���c�eJpt�T*�,���iϳ��`@�IǇ~8�&ΚU�z��.Q��/��1�2��չw`Ǖq̆9Ih������� /I	S�܊��\�l�I��0?�/���	H�aqe$�#��l ��N��dle�&3�����1�A���ckp��T�gt��c��4�p���1�����k���Ո%��GՏ������_�ͽ���8�jl@UU&���@&�Ғ�8�e��,��'�T����x�Pi\�d|_l<��gU�� a��nE(0D��k�fJ�z^�I�[fK��̶��N9�5�2�o .p�B]7}&J���Qݍ���ksL�3�]�{2��it^_���[���|�B��l(��!���B�������=��W��il%M��8Y����qC8Bk�Z`�H���ܶ�,f@Y6��q�<�8��f�=a|�H|پ�����.��^������I��Q[__E�����eEY�/#��$��S<?ɺ�Q��BAE!�tp[�e_]��>F_���+Z^^n�-#p�A��"�z�^�������5Ì{A�Z���+7��_�, �B�k ��Fvq݈�|{�޽�נ6�37w�Ὗ~z���z���ZO&��ɇ������-?|�������$>�<.`���X�ޫp�WZ� [�?�h?�ehO:4�#��?��c����x��ㄆ큍�[>Ӹ�2�������g�>�j���v烯>��'���LaK�N+���0 �Xݠ7t��G��mPzg:q�����qx:B�(5|��<_����ezcuz�cU���G?�W�~?n#���Ël �O?���_>!�^>��#��a/���ѣ�t�>���O~�˹}z�޽Ǽ�x¥�^��:�˿z��W4�d�G`#̆����K�;����I�!g��ˏ>���`?���h�_�+ؿ�W��ͺn�w��?������Y/k=h�E�1�)���}��`�����7 ���pN�;��������_�|���΅矟y![����W�?��'T:�V�    IEND�B`�PK
     ���Zq���W W /   images/7c9bed20-c7d7-43dc-b689-820375f46db8.png�PNG

   IHDR  �  r   5)�   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���{t��}������u�,K�,Y�K�6$�@�!�����4�%cH3�c�$�==s�G͜�4�9I�`;&�!mN��j�in��K�IHq�p3$˺��E�m����?d l,�'m�_k�%Y���1kyi���o�    �wy{�����B}.Kf��L���Um��To�jIU���^c��K3%%�L^#I.���0����r)/i���4��_�#2;t��O�u�h�ȥ���z0HC.�4���>�A��!�=��ߓl0;�9�,r��4�C2X[�����7��      ����+WU���+<_��bMII�BZ
fYM�P�e5&+X�5�� }���5~�ג̽���_��L��ߺ����rU���ܯ��
�^��_�:�[kX���ˍ>�Ҡ�!��d�2)5�I����on�|@���>I�if}I!�5����u,y�?X    ��b    e���\SSScP֤��(͒7e!4ɽ٤F���U/�,I��jcgOaC&fR�������i���������2;�I�-�,)�4wp$9�I������c��       �ޚ�V��$��4����nu.�s�!�2�u�LIu�>��je�)�L�kM�s�BG9��l@������}A��-y�{�ue=�vg
=-���(   [�  ���zݺƴ427UrJ4���� �u�)��Hj�݉�l��r����t��{�Bo��zf{<xo"ﵢw���ӱ�?v8      ��a^�����$�l��l�3�F3�-�F7�m�f�T+�L�f��I
��q�L�s�S��2uJ�ky�4�v��/Yf�z:n��c�   Sw   ��_S�/j~b�*��2͗Fo.�)NZ����}�>w�YP��vɽ�G���\}!�]�������Ñ�      �ym_�*f�s���T�z�T/��nj�L�f�����FN��4"�N�v��9���vȴC�vt�����۳ؑ   �d��   �N��k꫊vFf~�Kg���v�LgH����AIݒ:M�+��i��$Sg��d��ù���߸�@�P      �ܴ^���X��ZB��$���<�7K�d�l�ܚ}t�L�!�����&{:�=-Ϟ��t�7Wtǎ   &w   ���mkOJB�P���A�u�FOao���I;%�-�r�2e/ʭ+�l��v�;w}{�@�P       ��n��r�P�\�\�����[�B����u��I'I���
�}.=c�S�-X�M�=��q��y�8   `�1p  ��Ww������+���,;W��&-�dL3\zI�n�~-��z!1��S�U���Eݵ�;      x��6$IOk��TSx�����N�L'K:I�I�cg�ߥ'��qW�.��L���X�;v   p"�  `J��~M}����ȃ-�k��s�϶��2�OҎ#7��w�n���C�������     �i���5����[�|�曍���*�4I�q��Ϥ>���|�����oݽq�vN{  �T�   �V�u�GJ�E��"�](��}�X c/��)��_pٯ��7�*��М�ya[�ґȍ      ���6$��:�,���N5�i��ͤS]:U�<I�ȕ@Y:<zT����$���{:V��   8�   �.oϵ�n<�C�ăs2;0)uJ�&�w�iGRʶ�����~�^�     ���7��id�/��|�1_N`&�Nwm5�&ۜ&?������    �B   ��ᣫf&���`饞�e2] �2v���(�yw=mf�����?J�3���}Q��Y�@      ���ew�*M�H��p�3�~��ΐ��X/0U�$���2e�,}hw��=��   0�0p  ��hi[Ք)���/3�e��SR�����Y����s�BxƇ���+�c�     ���]���"�s<ՙ2;#Hg��t�ΐ4#v�q璞��!s{����{��;cG  ��1p  ��h��Wk�ʡ�%-q�ȴ@��	���H�M���-H�=���}�'�b�     L'uׯ�/}a�-��B�-��@Rk�6 ��i���ɥM�$ܿ�影�   P~  `l�mH��.3-1i���$bg���������k[�oWjۺ6�x^2�     0U���g��o��ۂ̵Ђ��6� �V�vH���&��������I   ����
  ���a��s�}ȥ��~� ��^���|��m�m�R��ӱrw�0     ��d^�W����������/�47v��6$�-�/����q�S��   051p  ��;|J{0��d���gJ ���ɷ�m[&�^SS��_�q(v     �xk\vGk��E.-r�E�Od�� $=/���;������o�  ���1   �P�GW�̗�t�Ur�+I�c7�1��]�c&L�+����;     �h��WkC��yJ�;�]��N�ΓT� �A��Mf��e��������A   ���  ොt������g�f�ߕT�	 �H��m&���[w�����۳�a      /=�=Y ��l�\�$�-)�n�1�I��K�V���x�3��   0�0p  �$�a�ꓓ,\-���t��$v L��r=������,�Gzf�'t��b�0     P�����'��J�p��_ �&�SRC�4 � n�[3���4�枍�;   �1p  �ƚ�V��Z7[&�"��! �lH��dz��	!<ҕ�~RK��a     `�rk�f��!I/ti��.t�I��� `�pm3�=r��]�\�   ���	  `����/�*T>왵���%�b7�1b��oq��P���}R��Y�0     0�4.��5��"���"3],�1v L!�]�[��{�߶+v   &w  �i��<4���p��_RE�& (\�j�G�푐�#]o�;
     L��mkOʅ���Å&]��cv ����#�}�S�b  `|1p  (c�׮���o��ZI�b� �4�W�Gd��+�I�Xz��o޺'v     ��jmR1�;R����Ã���� `���[��k���l�6  �w  �2Ӹ��$m.��2�#v @��i�f�oɤ�s���mKGbG    �7�|͚�����Z�E��-)� �]&�{y������  ����  �,l�P��h�n���$%��  o�d[M�c�~��?��X�;v     �]��k��.6��$�X�E��1`*�b�w�r`}����P�   ��   S�춵'�?��Ҥ�c�  NH����FOz���~䅯�8;
    ��ն!iɺ��r�H�K�Z,�lI!v �-; �z)�����b�   �a�  0մmH��烒-w�J�d ��a�&�G�m�����+�cG    0U5|t�̤��D��ʵ�LJ�� 0N\)غ�����o��  �c��  `�h�z���&�>)��= �(�2���l�+��{�O�    `�jX���|��>z:��2�+��W��-K�vu��|�   �9�   �\cۚ��[\�IIU�{  �J��~*�f�o��O����     �U�5k�{�ktоX҂�M �I%s����wm�eS�   �>�   �Q{{h�>������!�s ��HzԤ͒o�{Ŗ���;
    �1wӺ|c_��D�Xf���I��  S��Q��TUS��/|�ơ�9   x5�R   �HS��
v�I��uF� ���Jz���<<$���X�;v     �k�G�8��P��e�I~�d�$bw ��N��$I�]�,�  �Q�  &����sv1o�Iv��ٱ{  e̴C�˴YJ��q��     x���UMn�Œ]"i�K�K
��  ekX���e�gwu,�u�  �鎁;  @Ds��r�ґ��{Iu�{  �R�I���dY�e�ƕ�%��Q    �饩mu��]�Kv�K�� �(�������q���1   �   D�|͚�J�߹�&I��{  x��&=$�-�lsoǊ�1x    ���ew��'���D�Œ��_ &w�wC�g���'�c   �    �@�׮=W���5��t SC�\��f�@�9�W{{;
    0�4^{癉��\v�K�3���M  �M���=+7�  �.�  L��׮>'���\�KJb�  pJzإM��Ի��Q�    ��z�	�ҿ����M  ��-!���{���  (w�  �Q�5k�{N&��Ű P�z���L�ݵ��c��$��Q    ����A���$��	 �q�%s��ގ[�  P��  ���k�<3���d�İ 0�x����d��e��ގ[��]    {�V��s�_
���b� �fL�nB{�����  Pn�  �����5�i����)I��=  ��]&{P�[R�fNx   ����mu��]z���Œ�n `2p�w��O�l����-   傁;  �h�誙I1�'6:l��� ��e;%�ߥ�����]����E    ���Ҷ�)���u��+$��	 �I�(ٗ��>�}�'�b�   Lu�  N�M���}�n�ɚc�  0�vH�$��4���c�K��    `:j���k4\�IK$-q�|I!r  S�!�����u,�;  `�b�  �5��Y����\�c�  P&\���t��_̧����bG   @9�����bRxo��+l��%�bw P&�e���]=w���1   Sw  ��Դl��������-  ��Ԥ���އ*��?;
    ���I�z�e�%6zJ�bI���  (sO�§{6����!   S	w  �ct��w�.��/\�RR� �i�d�c�6I���n�X:;
    &��k��W�������f�n `�ڔ���y��'c�   L�  ��M���}�[��/%���  G��c�6�kS���G�ޞŎ   �X^3h����M  �����������Ď  ���  ���k�\i���tf�  ��H����OK���l\���A    0���>9��
3}@�+$��	  ��N�������u�<v  �d��  �(�h�ܐO?'��b�  ��ʻL��\���]�=�    NDK۪�4�.�%�ĥE��  �[�z(dي�o�;  `�a�  �J��yۜO���f��  cȴC�˴��������w�N   �7�����h��=��HZ����B�,  0v�&_���CO����1   �w  ��Z�־;�I��c�  �q璶��~��?<\|`߷>�/v   ����uեJ��Bz�g�~�I���  ��yW��g��ߋ  00p  �^}ۺ��e�Y���G  LW��?���٥V�qb   ��v���*�׆�Lv�ܮ��"I��]   ��YHo�]ۮ�!   11p  �Zӵk��k�I'�n  �Jj��%m��)�C[vv|z0v   �)�mCҨ�w�i�\��t�����  ����\�ձ�˒y�  �� �ii�G�8�PQ�9�n��  ���I�����`�g��p�(    �_�5k�+h�LK$-q�>v  �
�A���=+��]  0�� �i�y��\�V�I�[  ��5 �G.m������úky1v   ��^9hw�
I�c7 �)k����,����۳�1   ��;  �6��^;�����X�  Pv�%�ĥM��Ի��Q�p   ���ew��'����]W�tr�&  Pv�d���v��T�  ����  Ls��^-�$5�n  �B���i��6�v���d;
   ��kj[ݢ`���D�ߕ���M  `Z4�?��e�5 �r��  ����6T�7�n��  ���&=$�&)�AW�m��   plZ�V5�!wyp_,�%.] �g  ���W��7���mW�  ���/  �l5_��bw}]��[   ^�Ӥ�rm*&����W�;   �����3��Œ�HZ   LB�r���c�7c�   ��  ��u��}i�I&)��  �f\zҤL�`Z�����坱�   ��b^�W�a������z�L�bw  �����P�������  0�� ���x�g&�ΥE�[   N�Ӓ= �i���X�R�    �\�^���T�.5�.w��$�'�  `�2�0ˮ�Z�ñS   �
w  P6�,]{��_�4+v  ��4i�\���]�=;   �*Z�V5�%Kv��%.�/�  ���$�l���Ϩ�=�  p�� �)�����n��  0A��-˶��x��A   �d�|��9�g�b�~�x^  L�������Ov�  8<�  ���׮>'u� ���-   ј~%�.{�ݷ�v��T�$   `�4,[}r��e��R�]f�9��   ⱝ��u=+7�.  x�� �)kε�����H���  0�t��2m���9j�鶎�#��   ���|͚���Œ]"�bIb7  L2%�?۽��3jo�b�   /�  `�9톻+׸tc�  �)⠤��9S�`����ΎOƎ   ������E��K$�L�Hj��  0E�c���񉽱C   �w  0�4�Ѫy�\n��w�n  ��J&=&���lsa$���o޺'v   �zպ�be�����f�TR]�.  �)��Y�������!   Ǌ�;  �2���^���%5�n  (3�\O����m.����w���Q   (-m��\����er[,���   �̀�n�w�7b�   �  `Jhn[s���On  L�Nwm�i�ܷ��T?���n�  �)�mCҒu���l�4zB��s�s�   �tWw]r��Z^��  �Fx�  LjMm�g�W]�4v  �4W4��o��6[�?�}�'�bG  `�j��Wk�b蝲�1���+�!v  �4����z:V�  �z� �I��m�)%�ߖ��[   pT���ce�c�Qw���:����   ���k�:+���f�r�L�H
��   �j.�(��t��y�  ��a�  &��k�\��ߒ�9v   ��AIK�c7��H�����[�bG  `�5����$�BO�K2��fz��ٱ�   p�I����|+v  �k1p  �N�ҵKM�5IU�[   p�:ݵU��r�R��;;>=;
   ǡmCҒu���l���l��ߑT�� ��2����L!��f�p��LLvӚ4s��Us�2�X�����h_���{����!   ���  L"nMK���I�E��  P�J���i�e�5�m�]����۳�a   ո��$�\Z$�%��+�:v `zI�)I���`JB82NO��8=��瘤p��L��� ��Q{����e����fGF����R�*����Uʲ߼���,S���>0�\Z_S]u�_�q(v  ��p  L��pw����W$�h�   L�~I��|�����oݽ��m��   ����uu9�Γ�%r-6ӻ%͉� (fR.%IP.�W�����z���=��|��NTǨb)S1�T,�)��_�u���X�8-���#+��]�\�;  �{   ���UM��#�ݱ[   0i�ۿ��O%�txd��}��Ծ�Q   SY��>_�U�o�w��wL�H��bw ����M�$�'A��G�|?�>=��f)�I5\L5RL5t�-�w���<W�l����!  `zc�  �jn��mn�?J:3v   &�Nwm5�&m�\��ӱrw�(  �ɨᣫf&#�;��ȃ-�k���$%��  �K0S>��咠|��%ʽ�����z�d��0R�4\,ih$��HI�#%������U�ׯ�Q�  0}q�  DӸ�K�,��dͱ[   0euJ�f��n�J�u�ƕ�%�)Y  0m���g��s_3f?[���4̔��'����dt̞O�sA	�uHr������)ip����"���됙-�w�wb�  ��{)   ��ew~��p����[   Pv�Kz��[�����}R��Y�0  �ո��$�\Zd�.-�� v `�|��o��9q��J��[N[ǉ�2�P������h`�����t��le��+��  ��f  ���s��-��H��n  ��q@����gf��[x�nq��߿}8v  �Q]ޞkij9ӕ�'��]~�d�Kj�� ?fR>�9u��O��/<�t �,s��th�ݻ�    IDAT�������F8���d�W���)v  �^� �	5g��?����!   ����3A��\�P�'T
�wm\�d<=  &�춵'%�s��2;W�Εi��B�6 ��yy�^ȅߌ�_�>�=�0^�ԑf��������R^<��}�{A�J^!  L�e  `�4-]�g&�U�   �M4�i7mw׶ ��I���|�+v  ��?��ZU��/4��k����dͱ�  '�L�%��r��_�z��+w��PQ������{Y�{�g����c�  ����  L �9K���H���%   �[eR�K�M�Un�2���P�g���| v  �d.o�5Ϟs�_��"�-pi���%�n�)(	����_���Q;�Q���������e��w}����텯�8�  �7�  `|�mH���.����)   �8(�􌹞4�Sn�� =9�K�����Ď  �k^���UqV��r�9nv��Βt����} �c�S!��"�(��'A�|2:^��u�-K3׾C���?���R��	��U\���?9�  �/�  `�ܴ.߼����li�   `��|�L�ܵ#ȷ+�m]�u���v^� �)���5������m����Od?KR9 �&���8i�ho��0�ճP��N���i�W������!  �<q  ���n��rp`��]�P�   `��7�)7=e�oϤ����j���g�;�� ��������tN��� ���96��>v ����������|�p�:0�����?���!�Ǯ��ʆ�+TΔɶ&I����Y��	  ��  `̝v�ݕ���L��   �BRI/��K7=�rNY�\�l{Aw-/� `�kې�${Nv�oW��fo���n:Ǥ�%�c' ~[L�|��\�B>yՠ�"�(	L��h�����C�)ĳ��C��\�BU����\.� #w  0ָ�  ��¶�n�n4��n   ʉI}.m�i��vȴ�3�H�<�ױ|�>  &��m
�Y�<%�/�|��K�7�ΑT9 �
I0�s��i�Gy�O��ePֆFRu��ׁ���)x^T64�0#w  0��  ��v    ��$�8r;<�W�]�u����,r"  c���5����[���b��:MR�� �����$(�U�GOa/��s��`�����ۯ�b;�#�//��I���Y��\�,a�  �
w  0&N�rU����>�}0v   �W9$�s2�0��]��.�hn/fI�W�g���  0�4��nI�Nβ0ϔ���N1��=���f�n H�L�\���[N_p<ܥ�}�Գ@�k�j���G��<���T�Kf?��%/}��=q�  @9�$  8a�6z��C҇c�    8nEI�&풴C��L�K��i����w�����2 `L�v�ݕ�[�h������#'�K��N�4#r& @����_q�zE>Q����\��|;@�.���9�}�҈���G�MF�  `�1p  '�u��}�F����   `��K����^���,�Up������������"7 &��n��r�P��,I�Y�S]:�d���3;���\���	 �S!��"��p��z� �'�\/���ރC�S ): /���?GF��g##C���O훸:  Pn�7
  ޺��д}�7LZ;   @tC��Lڕ�:-h��;�՗ۥ�;Cf��f'/���ر ��3��UŬrn�U���[e6�M���>������-��' �4��|N�|�B.(����|d��`
�=0�]{�弶\Ti��or�~R��z����˗�t�쟘:  Pn��
  �"�9K׬�ly�    S�I}.u�� ^��L���;�m��Yg)�}��o플��`��v�ݕ�C�J���y���y�I����Ms�:YR>v/ ��^>����Se>9<fOT�O8�@��,ꅮ�J3&��Ӣ��=���GF��f�?���o�:  P��7  ޒ9K�~N�?��   ����k�I{M��f{\��2��=A�׃�����|޳[-{ձ�M���s��w�	����fg�}�)kp�l�$k��l3�vi��FI3bw �]0Se!���÷ÃvF� �������ܯb��N�v��C�������T���d���Z�  ǋ{�  �5/]�����    �:�IꕴW�=2�k�W���{C�=�|o�'-%�ܭߒ�A^6@l�W��Ns�����>ە5��l�7��`�l�7H6[R�F�<� e�c�ꊜ*�9��憋��۵���K�J��q}���}�L��kÊ��*}  �xp�  �9׮�En�cw    �8��'Ӡ|�}w�Ӡ��̽ϥ>s�I6����՗��\6�˲�R������mK��_ SҼ�/T�WV泴*W��4X}0�gf�&��L�n�7Y��UnV���ToR�KU��5:T���� ���OTS�WMe�1; ����T�u�S����I��%?�?o�U)T�����w�m�  �w� �1kn[s���.)�n   �)����2;$WѤ�L�L�/I&�IRf:`R*�C&q������((�^��,�3�\!;����>��l8ͧCŐ�6`�������3�(Kuׯ���
E��U��,�,�*	�d�,IrY��I3B���U�Y��*�T���j�f&�W�LA���.U�T)W����7  �[!����pd�^��; ��ᒞ۵O�s(���lt��Y�Z�r�L��]n��ǰ  �1�  ���,]��L���
�[     'lĤCG�����[�xwi`��P��U������f�Q��p�Rz�� `
	f��̫�����U��I 0������bg�=�J�������Z�B��tcφ[�f��  @c�  �T�5w.�$<�/�        �De!�����TU��xv ��K{�ջ��^�c�Ӣ��='�}Be�,_U���+��� �2�]h  �������ǒN��       �de&ͨ,pJ; L�,s=�R���i씲5VwI
U�d�ʃ�}=�W<:&�  �%�  �u5|t��\1���w�n       `�yy�^7�Bu��;	 ���ᢞݵO�Kʓg%e�z�軙BU�,W�LJ�{:��Wc� @�a�  ��u�9�Jߕ�wc�        0�̨�k֌JF� 0I���מ��3����%)(�4H!�d������1��  �LpO  ՜��W�       0�"����Fg�ܠ�ϝ�ٵ���`�h��V8�s<ؘ���)�yvN�F�[ض�0�   e ;   L>MK���\��       @LI0��V�~F��+�s  �#�5�U��o vJ��q��\�*�SR�𾞰g����"  `*Kb  �ɥi�>h�/�Wz       LSU9�4�蔦Z��T(��u ��*9�90$�Rn��#����z&OK
��w�X����}�'c  0U��<  ����/-�,�����[        �H�FOko��Tu/� Sѯ{���P쌲���H�����|�B�����������  �)��;  �$�^������5?v        %�j�Y��3���B��l`��g^�;�줇�HYqܾ��)+T4��vݻ�q�  �2B�   0	ܴ.����3n       LU9��T�sN��9���@���+�c5�l|�L����p���CK۪�q�  ���  h���.���       ��V[U�魳t�I�j����k��RWS;��XH����~yVz[j�{uy{n�/  &5�  LsMmko���;        O�U�q�,͟[���|� �8��*�N(?�|���L�@�̳�ϙ��_'��  `�^  &��k�\,��3       �L��T��晚3�Z��@�K��g�`��⩼4<��%�|�{j���Cۿ��	�(  ��x�5  ��9�}�Yi����n       `��V��P��
Nk���/��p1��Q6<-*�3a׳�������{W<1a  ��D�~  �l.o�YZ��q;       ��TW�����4n�v ���
��	e��ľ���ˋC5.���m]݄^  L
�4 �44gN�_����        ��B>QkC��j*b�  "��8�sLY�y6a�̆�+��|����#���]  D7���  D7g随H�ג,v        '*����F�4ժ��3�  �p)�����e�KÒ�|��|�Y�64����'��   *�m  L#M�|�K���jc�        p�f�Th��*pR/ ��֯���(+��yq`�/�T(��O3�z;ny`�  @�� `�8��U��z1n       Lq���No��S�g2n ��$p��X�$��鰲�CI0}���u�q"  �D�>  �����J~A�        ު`����yR�j*#�  �^0�c.��]���FN*�ҿ����  LI�   0���|���Zw�       SҌ����R���
�[ ��R�i����e�,�G$y��{:�P�:cƹ��?��{?�  &'� P��hռ`�1n       LA�L�j����T��7 ��K�8#첗��]�S�����5_���x!  `"0p ��]ޞ��r�H�; ����;��,����;�n��K/3==��R\d-�,QR$[�I۲�CJP,[�DQrl�p;�3�_�9�a�A����ț ��+��Erv���޵޺�9'/zHΐ�TwW���{�h�@�C9Uu�{   �v�tZ��=˱:?�:�1p?Y��6��G��mUU�O��YL 'w c뛛OFď��     �ۑe�Wf�3��p�܏G�{DT�ݨ���Y�[ ��c� cj�3O�����     p;ڭF<tf96�f"�R� PG��0u�X���	QlEV���x��_N� w C����g�����p�    ��X���#g�c��L�@��E��e��ܫ"ʃ툪z�̅gΥ� ���; ���?����Sw     �adYęչ8�����v �N��c�5;�""�D5�.��œO������ ��槟�dVů��     ��h5�x��r�/N�N`���ckT���NT��'7����S�  G�� �ș�>�VE��Sw     �a�N�⑳�1�i�N`L�t���Z�hEd�29+��nE����|���S�  GgT��  ���(���S�;     ��,�OŃ�����kk ���~/u����s�=�A���NUV��/|��: 8� ��X����BD���;     ���Z��s��e�K '�A��Aꌱ�5Gh�U7�r��+ٕ��� 8 �X��ԩ<˞�"�S�     ��ɳ,�m����h� ������3�_UF�{9u��e�ḫ˼������}� ��� c ��)�v     FY#��Ӌ�� ������A�ɐ��vꊷ��({;ͼ��i��3��9 ��1p��[��ӟ�,~!u     ��V#�N/�씽 �����eꌉ�5G�k�`?�����7ʿ�� �;Y�  �Ν�s_\���Dd��[     ���[�x��btZ��) �������z=ʪJ�29�"��+�+�Wֈ��Z/����x�sϥ� �� Pc�v���    U�V#:�d����������7"��߫*���vʬ�'�䓶q PS��@M�?񥟍*~%u     ��v��^�Vӯ�8>�vb{��:c"�ͩ�	���EU~d����L� ܙ,u  p��>�{��T�?FĹ�-     �ݾ5no�p���a<���(J�ۓ��(v�D���?kDcvm���_�7^I� �O ����ޓa�    �j5�x�Ԣq; �jX��ҥm����<��N]�Ϊ"����0+�a� ��y�  5���ӏG9u     |�f#�O/E��H��+�*^���A�:e�孩�	���GU��槟�d� ���@�TYT�#���     �*ϲ��Ԃq; Ǫ,�x��V�R�Y�Y�wQEy�Ud_����?�� 8<w ���O��_�"~<u     �U�Eܷ�3�Y 8>ߺܾ�5nY���}D����se�o�N oT?> |�{.���~��jD��n    ��:�6kө3 c�a/^ڊno�:��R{Qvo��xy4�V��<����[�� x.�@M�����     �����v ��~o_�q��ʚ����:�=�Q춋*�݈�AX ��Q�� x��_�������<�f�G#Ͼ�����Y    �6sӭ�w}!2O�8&W������(J�'iUQ�SW��rY�u���������?H� �7� `�=�d���ƿ��L�^�e1�n�T��V#��<��F��y�y���h7�h6�h�ydYD����������UTQEQT�����3��c0,�7(bX�'��   �I�j�����h6�8��7��ͫ;��?£i��,�ػ�����ḫ\��G�����v� ��5S  �m�+��Yd��0�ڭF�M�b�ӌ���?S�fLw��i�˒n��h��_bn���������� �{����c�7���A���   �ۗgY��\4n�X\�9����𩓼��D��%�F��n6���""�v� �ݹ� #l��SsY��QD�I����g1;Պ��v�O�cn����h5��˻��b�`7w{��ߋ�=�w    ��=��:?�:�1�����vc�`�:�;P���L��>�ḫ���co���|)u ��\p��g�ߪ���DeY��T+g;�<73혝z���u�ȳX�i��L;"�#�ֵ���^�����^/���QVU�P    F��lǸ�#��q��^\�9H��]Ț���Q�S�Ceow*��^D<�� xg.���ڼ���s�p�y�3�X����ܭQ�8\f?JeY�ͽ^\�����.�   L�V#�G�Y�f�34 �^Xƕ����}��Θ({�Q�wSg��|f5����+_���� �^� 0�6>����/��q4�i���L�/N��\'�̷ŷ��ƕ�ݸ��7w{8   L�N/��t;u 5w�/���~��=�f3U��y+3����� �|�L� ��% ���O?��DT�&|��#�l䱺0��ӱ�8�V#u��e\���_��   `̭-N��չ� ��N�W�����O��1*�7���x_��bDk�׮|�7�i� ��� `�T�槟�wU��S�@��[��\����X��J�3z�".^ߋ7���N׃i   �q�n5�ѳˑ�~����˸�s�w�?(R�p�������/ˣ1�~1������7�R�  ��L  ��槿��*2�v��fK3qjy6V��OZ�Ո�q~s!�q��^�vm��j   �1p�ڜq; �V�Ul�����A�v�s8aY���"��k_�Q�wO7��߉��6u ��@ �(��gZ7��"��)P��wF�F����tc?^��7�z�s    �K���os!u #nX���ߏ�^�t�QU��H�t�<�J�qY4fWw���Х���S�  ��� #d�F����a,̴㞵�8�2��FV�eqje6N����~?^��o\ߋ��T   ��,�ӫs�3 AU��c�ۏ�� v�����5�ۉ���)��7�M-�͈���5 �-�@ 0"�/<5�e��#�T�U�F�W�➵���j�����E�vu7^���A�:   ��pfu.��Sg 0"z�"v��ߏ�n�A�S�ۍ���:�P���~#ڏ]���!u ��; ��,��zDe��`i�������Ld��h�]�و�O-�}��՝x�Ҷ�;   �j���`�0����no��A����0�A1�׸%yk:��^D��!��^��i���R�  .��H8��gֆE�|D,�n�Q�ek�q���X����UU�_ۋ�/ތ��;   ��8���s��L������3f���q���b�ݭ������O���h}�ʳ����n�I�; ������̸"��gqje6��X�٩V�N@�eqvm.ά��   ���vӸ`UUDoP��`�~�a�E��E���_�<7�    IDAT٦~��lm�eo'oή���S� ��s� [��?:����#b*u��n5⾍��gm>��<u	�e/_ގ�؊��0    ��O-��L;u w`X���1������c0,S�1����E?uơ�SK�Ο���o���[ `��� ��U�o�q;������b�[��<��K"�<��O-ƙչx���x��n8   prf�Z�� #�,��U��m�6f�����۳Qv�1p/{;�hN������[ `�Y@B+�y��f�}="�畉�j�qn}!��\��a;�ag�_������K�   08���� ǡ,�(�*��֟���(�w��o�{�)uV�]�(�3%�Z��L�ؕ���� &�� �P���V�3aZ�<��\�s����L;��#���{��nDoP�N   [S�q;0V�5/�����[���u@^|���|�q�w�΋��*�����?��n��:��$��3Ql��8������߉��I� �ʢ 9s�sì�Z�3!y�6���B4y�j�(���k7�WvR�    ��{��ce~*u�����uɼ��E��ͫ�e��ۮ����[����ؽQ�㐑+� ��� ��0���̸����8�޻�m�~rwy�ݻ��g�W���A=^e	   P�F�s������9N��7�g�a�a���X�-��=U�G�n]q����ө[ `�� 	�y����=�����v<z�J,��,G�,�x���x��׺   ��+���4�:3U���������[#v�xaBT�+�Q�.9���ў��+_���� &�� ��0/�����_�f�Z�s�Scy���g����\|�嫱��O�   P[y��ʼ������h�[�ް������ ""�<��tT���%�R���њ���n�I�; ���O�md��z;c(�"�m,ă�����V��SUU|�������)    ��4ۉ�6Rg #lX���o���"E�C؁ë�(v�DD=�Ƒw"k�����~�ߦn�I�; ��FV�NDf��ؙ�n��[������eY��]��������FP�N   ��e�ہ�����������K���%v�dyd�����%�R���ў���[ `�8�	 'h񗾴���1���J�eq��Ÿ��Bd�o/I�?,�?�t-�m���(   @j�F��[��`rTխg��A�a������'�*�Q�]M�qh��b��;z�_��WR� ��p� NPg��vDe���X���έ��T+u
|[�و�=��\މ��v�/c    ���\Ǹ��;���8���dy3�щ(z�S���f���_����� &�� pB�|��t�RD��n���l�����gm.u
������/^�ޠH�   0��g9��n�A��2�Et��[\dFXU��ܿ�:���A�9������+�[ `xJ 'd0S�ZV�S���x��Z�t|+��[���}����^�[{��   p�ڭ�q;��`X~{ľ������C@�d�vD�Q�S�J��k[�5"�Z� �.��I�ē͍���G���)p��,⾍�x��r��mUU�s�\�ׯ�N   )k��qv՛aTUU��"{�7���0Jgف1P���L�qh���~kj����߸�� Ɲ���	����L�ScS�f|��Z,�uR��ɲ,>x�j�O��k�]�J^   �7-�x����"z�"�{��ڍفq�5�"�fD9L�r(�`ofؚ����oR� ��s� N�慧�]�e?������L|��j4y�8W���/^�aQ�N   H��g����"�[c8qUq0�5`�w��`ՠ��V�C˧W�v�o>�׺�[ `��� ���g��DYV���N#���V���l�8Rk�񃏞���rt{��   p����pB���W��{��;DQ�d����NDU��D�`m�X������- 0�����e�WR7��j7�#���L;u
�٩V�ࣧ���r�t��s    ����GUEt���;�Θ}0��p��e��f���9�jxU9�;�?��|R	 �����1:���ϗe���h�n��Z[���_�f#O��nX����_�����)    '���]�N��k�[�a{o������2y8���b�jD���@Yk&�ş���o��[ `\�� Ǩ(����S#�7��˩3��4y��Û�^��o��   81�Fn�w�7(b���A{o�a�$�z���ZSQ��jЍ�3�W#�� ��� pL�>�{��T�ՈXL�������Vc}i&u
$��+�⵫�x�%   ��Z����ͅ�0�*���y�}����0P+e��Ո��+0��|��Ǯ>��?J� ��w 8&��ޯU�q;�o�ӌ�>��S��)��έF���˗�S�    ;�᝕e��a��c�;�noeU��%@��ȚSQ��K���g����#⯤n�q�; �'��7���ZD<�:���l'>��z��^E���oƋol��    8V�]����;|�B�n�֠}�``��HU�ܿ�:�����as����_,�s� ���n�\�q;#mci&>t~-��g�:�a�   ��,��n�3��*b�wk�n�0Z�F+�ю(��S���ϵ�S��0u �w 8eY�Ff3�;���޳�:F�Cg����x��v�   �#�n6�3l&IoP��� v�����GQ����=e��(Q��ET_��|q�#� ���<uo��^��F��nY��=+q��|�����z=^���:   �H-�v���B�86â�݃A�9h��I ܆b�jD9L�q(Ys*bj�W������ Ɖ� p�e��a��ʳ,>|�Z�/ͤN����{W""��  ���iy��x�����A�toڻ�z�"xgyk&�^=޲[{�W��"�� ��� p�>�dscc��8�:ު�g���cma:u
��W^��_�M�   p$�]������pW�E���o_i/�*u G���ػQ����~3���ҿ��˩S `\�� Gh}}�φq;#��g�7��
���[�aQ����S    ��T�w��_��~/����w0H��qɲ�Z3Q�kr|��m�ss1"�^� y�  'Y�K� o�j���7���|��Z,�vRg    ܵN�4�,����ūWv⹗��}�z\��g�0��LDd�3�*"��'����#�* ��'�y0��'Sw���y|���X4ȅ#���6�٩V�   �;�gY4�ŘHEY�ͽ^�re'���x��v\�9�AQ�N�$eyd����7����� 0.|4 �JU|.j�r�]�Ոxx��X���Gڈ��ވ��H�   pۚM7�=â���~l��b�ۏ�J]�(��3Q��3�D���G���� Ɓ �O<����x5"N�N�V#��?��3��)0�v����R]�   jf�ӊ��.�΀˸�׋��^�R� 0���ke=�Nd�a֞��ʳ��F� �;��#����sa��h6���q;���v<~~-2   j��;	e�w��7��_��_�5n�=���	�V��,�_J� ��� 8U1u4�,>��z,�ÉX_��O�v   �K��WĜ�������+Wv⹗�ūWvb{�U���:�ZSYM���(��_K� ���A �Kg��W�����*&�<���\�����)0q��ū�ƍ��    �rjy66��s	������v7��zQ��� ܹ��U���ɚSSK?p����?�[ �Κ� ����W�2n'�,����k����[��� ����S    �W����񩪈��^\�>����e ��5EM�հ�j�"�� �BM�� ����WS70�>x�Zl,����y~`=ZM?^   �/�o��eW���\��/m�p��ƭ��PE9�}����B'u	 ԙ ܅�'�������L�O/����0�������1   0�2�/8BeY����^�ׯ�Ơ(S'0��V}�f]{�[�O�� �:3p��Ш�_M���:�:�^L��ii��YJ�   �|@��rs�_����x}/��� ��َ��3�D�)u ԙ�; ܩ_�UE|6u�ii�8��:�.�7b}�>D   ��c������k�݈�/m�`h��I��v����/<u*u ԕ�; ܡ���D�Z�&��T+>���W	È��}k�i��   0q\p�Ne�^ى�/ތno�:�	��j��mD��; �����Y�z;'����#nD���8U�f��54    �ƍ�^|���q}� u
 �,oD4ک+�*�v9u ԕe ܁��Ϧ"�O��`��Y}p#f:��)��X���N-��    �eU�N�F�E/]ڎW.oǰ(S� @���ǰ���/<�P� �#w �{������L�G�Y���N���8�+�S�3    ަ,�9��n?������K� ߖ��"�zLުa/�j��� p��� FL�B9QgV�������mz��Z�~�   F����x}/^��W�9Ydͺ��~9u ԑ� ܦ�_��BD���L���v<v�J��tZ�x�  ��;�?,��ߌ�7�S� ���Zө�����>�� ��� nSc��ň��G©�V#��p=�<K�ܡ�+���4�:    "\p���t��o^��� u
 ���ъț�3��E\q��e� �)�곩�Y���k1ݮ���]=vn%Z?~   �.���lu��7�����Ț��IW{�Q�h ��� né_X��O��`2�j1���z=�ݵ����{WRg    DP�N`�TU�k�v��k��? u���3p���{6�x��Rw @���m��柉�9v3�x��R���Z������   ����󦢬�K[qu��: n[�7#�V��)�Q>u ԉ�; ܆�
?tr�y�=up>pn5ZM?�   ��e�F@oP��_�����) pǲf'u¡�E�B� ��
 8���,F�O��`�}߽+1�� G�f��]N�   L�����'�~o�x��k� �^֚J�ph��ྍ'~��Sw @]��!����N��x�X��3�s�3�ctfu.�����   ?��a���⅋[1,|�����fD�J�q8� �����3 �.����|� �[�Ո�[M�����]�,K]   L���'��^/^x�fe�: �Lͮ�� �!��!���33�3�;o��_�Vӷg0	f�Zq��B�   `B�R'p�n������Qٶ0f�f��E���_z4u ԁ �`�����I���:�6+��y�ܽ��,E��H�   L ��ru���0��FD�L]q8E?�j�; ��; F��:���n5⑳˩3���3��   ���e�N�������� p��f'u¡UÞ�; ��; ��^�r;��������]�f÷e0�N��z{   ��+���ҍ�x��^� 8vY�>�(]��/ܓ: F�% ���������������X�I�$��=+�e�+   �Ic�>ޮlu���Y�u��U�^�l6�t� u��� 	�?�����l��ع��@bsӭ8�2�:   �0;]�que��_�M� '(���NqHU���O�� �Qg� �#��9�]�N��:�Y�F�;   pr��8��38b�� L���I�px��'�|�����`� �a��*N���Y���=k.6�tZ�8���:   �0[{��	!�v &Y֨���j؟�w?�� F��; ��<��t��ӣ���N F�����   �	�i�>6���xy#"o��8�2��}*u �2w xUT?����sfu.f�sA 8�<��7Sg    �?��~�:��t}��� ""k��w��p��U�� F��; ���_��B�;/�<���,�� FԽ�s1ө�u   `l��^k7v{�ͫ;�3 `$d��ܣ�����J� ��� �Ec��Saeȑ���btZ����ʲ,8�;   pr�mw��RWp'��z��m� �MY�F��/���I� ��� �E�ϥn`�L��q��B�`ĝ^�u�   81��������nw�\�1n����>�c)��ϧn �Qe� �*�����G�.G�g�3�����    '���~�n�~o/���u; |�z]q/?�|����w`� �`����I���X�����L��&ά��t��:   ���0��38���0^�h� �&k�S'Z5�7[1��� 0����T�O�N`�<xz)uP3�o:�   ��+[��	��n/��Ei� �Q�Be���Ϧ� �Qd� 2w���l'V�Rg 5sv�w   ��l��\qa�A/^܊aQ�N����͈�F��r�S� `��9 ��^�r;�������κ�ܙ�   '��k{�x�a�_��v 8�����Ъr���t� 5� �]�Ƶ���������X�s��3gWg��j��    &�~o7v{�3x�aQ�o�`h� ��5�3p�r�p�'Sg ��1p�?�:����i�ہ;�eYܻ>�:   � ��FYV�3�[���/nEoP�N�Z���	��,����w�2w����t,�uRg 5w��|4�,u   0!�2�luSgL�aQ�ol�A�: �'���=��'��� ��� �����j�����N-�N �@����չ�   ��ts/����e/��ݞ� p'���9T��S����� �Qb� o�of?�>rg;��G澍����   ����x��v�e�:e�e/\܊�� u
 �XV�+�UE��gRg �(1�������������12�i���t�   `��E\���:c��e/�a� G!���="�b��� 0J��-�*7p�Mw���4�:3�6|p   8YW�����ΘEY�ol�ށq; �F��Q?�x�f� p|��M�\�'+�SwP�֍P���2?����   ��y��N�eꌱV�U�pѸ �R�5R'ܖ�̞Z_�X� � �~���𵑻�j�qvm.u0���   8i���.ތ��R���aQ��o�~ϸ �T^��{DŠ�S�+ `T�����O�@��]��F��� �ԙU�   N^oP�K����q?R�a�_܊no�: �NV��{DY>�� F��; �)�ܹ;Yqnc!u0�y�˳�3   �	��īWwRg��ޠ�o\�}�v 8Yu��eU�#q���[��1��Wq 8&��Y�,>���z[[��N���x�]�K�    L�;�ƍ��������oFP�N��V�+�U1�_o\�[ �0p���h�埈�z�t��9�6�:� Ks���n��    &ԥ��ڵ����w0�.nŠ(S� ���j6p�(#���T�
 � UT?���zk���8�:�g\q   ��ՍW��DU�.��k;��ś14n����oW�?�� FA����q��M�@�ݳfl
��3+s�gY�   `���9��/o�BUE\�����  8Y5�W���#*�`���8 ��~���죩;��,sM8Y�fK3�3   �	��׋��r��=e/]ڊ�7�S� ���j8p�r����?~ u �Vï� p�v���������tL���3�	sj��   Ho�ۏ��v#�{��)#�7(��ߌ��~� �Ly�qUU���x5�* G�*㏧n��κ�$��8���   ���2���MW��bk��x�f�S `r��{DTÁ�; ��_��(eُ�N����<��Sg (˲X_r�   Uq��^�ti;��J��LUE�vm7^��âL� ����j�é  �z~���C����t�y�:�P�WfS'    ���^/����q}� uʉ������o�խn�  "��ܣ*[��׈0�j�U �ƙφ��}    IDAT����I�A}m��$�2?�V#u   ���2^��/���A�:��UUĥ����nD�7L� |[M���F��� ����hE$u��l䱶8�:�p�ˮ�   �i{��������(�*uα���k�݈7n�E5�������#������ �R3u  �T���d�8s���#��C`<�^��W.o��    xGUqe��wbmq:�g�����jX���qs��: xOyD��#n[�c} L4w &ZVV?\׷������(X�i�T�}��   FWQVq��~\�����T�-�D�Y���2.�܏k�]���,��_���R' @J�{b  G�ןiEߟ:�zj5�X[�J���(   PEYŕ�n|��k�ҥ�����b(��ڵ���W���-�v �����r�z�3O�O� �����Z�.�e����td����hX_��W���    8��������^/Z�<��:�8ۉ٩V괷������Al������SQt0"^J� )�0����g�ܩ�ג�ѱ2߉f#�aQ�N   �m���+[ݸ�ՍV#���v�ϴcn����_]��ck�7vb0�� H�*?_N� )�0��*>���zʲ�����ёeY�.Lť��S    �ʠ(���A\�9����v3f:͘�j�t�S�F��Ѿ]�7(b�7��n?v��1pD  �G���]6 L,w &V���(KB3�h7�3 �f}q��   ;�a���GD��yL���j��n6��̣�g�l��Y�o��,�*"�����"�����������^��n�x �H���G"�,"�rz &��; ��ןie7��Π���S' |����Ȳ��#N   `��e��� @-���]Y,m^���K�Ƌ�S ��  �����J�A=�.��0z��<g;�3      8U��J] )�0���x��e@
�0o�      ��,�����(�X� H����TUa��Y[4F�ʼ7L      |KUU��NU�6 0���TK@=-���kq����      �AUUN�  )X> 0y.|���Π���:� ޓ�O     ��r����M� '�����W�����O����T+u�{Z��N�      0"��w�*#�|4u �4w &N��WxqG\E�`ua*u      G�����8� L���>���z2p�`v��V#u      G �
 &��; ���]p�,����:�;     @TUꂻW���N ��f����]p��eY�⌁;PKs�      c0p�x衟��_V0Q��(k�����������L'�<K�p(K�8     0ܫack&>�: N��; %��+en��L;u���M�����     0��`�1��h� 8I L���p��i~����     &�8\p���[ &��; ���>�:�z��j�N �-K���	      ����=�����b��D���`��in����E�    �I6&��#"���R' �I2p`�dY|_��g�ӌf÷M@�,ι�     L���WUqj�S�7�� N�� c������8������r���v�ӝf�     �$���dI�����{j�@��,���n��
_Co}����+_����޵7��>��Z�@�#Hb P�5�|��>/(ɢMR@!3��/�'��!��"DdU�?ߓs*�0?�o�+� lw 6Ƶk�\o�J���W:�J^��     ��j�G��t��� �,� l����;Wr뺁(������/     `C�\�`���w���a����ڊ��n`=ݼ�S:�Jn]�-�      PFm�G� �� l����q%7܁5u��     �fʕ�sJ[� �������63W���;�~d�Ӎ��     �)��s�s�Q��/\g`#X: ��ۿ�����t��ƞ���v��n�     ���{i��^�{ `#��^9��D��O���v��gr��^�     ��l����?/�  �`��F��iV���t��E ��yw     `�
�]��c� Xw 6B��ߔn`=����[�}Q     �@�/]0wMJ?-�  �`���h~R���tso�t�3�q͟c     ����{���� �� l�l�Ε\3p�ܵ����jJg      ,ON�KW�]��K7 �2��ܹ��?.��w     `��
���ѷ����^� X4�- ���؉�+��z������n^�-�      �<�ҁ{�M���t ,�� �{����ADX��Ԛ&b����M�    �M������oJ7 ��Yl����.`=��l�N ��.�     $�z�� ������-w�doǏJ@\p     6J��s�Z� �j��5���+����P��     ��)�NX�&7?*�  �f��hܹ�����	 sq}ןg     ����{?,�  �f�@�r��t��w�M�Į?�     �M���G��N �E�p �~M��t�iJ �ϵ=W�    ��SD������o�ӿ�Z: ������_�����F��Ӗ�;P�k�;�      .�|�=""rL��?*] �d�@�vg���\�֖�;P�k�.�      u�n���P5w �����n`}�����     ��_p�H9��t ,��; Uk"}�t�����ގ�;     �6`�)�B P5w ��#\p�ʶ��T����;     P����	�4����mP�&·�y.������     �r��s��-�  �d� @�w�l�1p�k�     �.����]�)�  �d� @岁;W�#�N ��mw     �r9��=""r~������ �E�p �^���VD�Q:����ہ���     T/u��$mN?v��jY8 P�W��oF�o,se�����_�     ����G��~P� ���z���N`�ٷ���jJ'      ,L�7gྵ�|�t ,��; ��N��K7��rX�u���+      P����޿Q� ź�z����g���;P�]w     �V9G�t��䰉 �Z� T+G|�t�ͼ���VS:     `!�]o��h"�D P-w ����2��w�6[��;     P����� �2p�^�1p癤l�Tƾ     ���]p���� �(� ԫ��<��7p��;     P��o��=7��� �(� T+G��L�>�N ����     �UjK,U��7~�_���� �� T*7MxϦ7p*�e�     �(����,��� �E0p�Jo���x%"�Jw�޺�qo� �۲p     *���tByk��� �� T�O�[�X]�K' �U�     @}rjK'��$w �d�@�R�^:����.�ui��    �m��H���	 �� T)5�j��_�܁�d�      *���S��J7 �"�P��I�<��#�d
�#Y�     ��9"m��&�R: ���:�������}���1p     j����?�]p�J� T��-e�df�T$y*     P��o��=7� T���*��w�c�����T:     `���tA19��� �� �)��;s1u��Hk�     T&���	�dw �d�@�\pgN\pj�u�     @Er�ț��n��; U2p�NM~�tup��E�9�d�     �#�]�Ҟ��?���# `���Sܙ���;P�I�GΥ+      �'��tBq����� 0o� T��N~�tu�u�u��|a     �K�f���ى�J7 ���P�q�x�t��6��v@%��H     ���h������P��ԿX��z��>Rʥ3 ��x�^     �9u��s�m$ ���; �I��~yc�\qj0���     �H�ODDΎ Pw ����F��b��`4�&/     P���J'���F���P������\�����N�    �z����s�� 0o� T'�-��b�&.�kn2��R�     ���)"��+V��� `���N�p����k�b4-�      07�s��O�H6 T����lm���O܁�v>4p     �{�?I9�H Pw ��s�b��b�����7y    �z�-��J^(  �f�@��Nf��>Ŵ�Kg \��;     P��#����4.�P!w ꓳ���p�`='mt}*�     0��Qn��K7 ���P��㷘��؛$�z:NK'      �M�=�������; ���7�n85p���ț�     @=ܿ�i�f� �7w ���s���`�M`=�\�K'      �I����%���_�P/l �����N\p��p��x�M^     ���""��X5�kp����P#w��R̺�t�S9v�     �H�=y�����K7 �<�P#�Lf!cW܁�r|n�     �#w��	+��M�J7 �<�P�����ۥ;����5 `}���l�M^     �9G�}���.�Pw �2�u������X#'�H9��      ����"�g_�I[� T�������~ica�G.!���b\:     `nr��گ���	 0O� T�iw�Y�񴋮O�3 ��ѹ�;     P�ܷ�V�V�Pw ���7K7P���t�_ur1�Yۗ�      ���"���W�� �����4͖�,���c�շ:(�      07��9��I�7p�*� T�I��,���w`�����|\:     `nr�sگ��� ���; ��7JP��7N��vp6��O�3      �&�>��:M�� `���J�f�tu�̺���� _��ɠt     ����Ed��~��V���P�&ǵ���l0)� �m��     T$w��	+/7�����P�&�_�X��Co� �i�t9��      ����J'��&�� U1p�*9����¹���ώ/K'      �Q����+/���Pw ��le���p�qm�Jg |���(�Ӯt     ��䮍���5Mv����P���_�X
W܁Us���v     �.���NXM�N �y2p�*M4�,���t��'m<���     �.�����
O��*� T%��,�!)�J�\�N      ���G��t�zHa+@U����,��x]�Jg Dۥxt:,�     0W���'�� ���; UI�[,G�'�P����2RΥ3      �*w��	k��.�Pw ��;�t|1.� l��r�;�,�     0_9E�m銵��q���P�&�N`s��}v<�Yۗ�      ��ϯ�{���y�t ̓�; U��k�3k��] ��9ǝ���      s����'�4[M� �'#@ ���kK�;Pʽ�˘��     T'G�f�#֌� u��@Ur�嵍�2pJH)ǝ���      s��6"R�uc+@U��P��[�,��`}ʥ3�s��2f��     �ݤt���ۥ `�� ���6�*�W܁%J)��C��    �:�nZ:a�8@e��P��k�wx6*� l��    �Z徍�>yZM�4� `�� �J�^�X���q�Kg ��R�yt^:     `!\o�"[	 *���l��n�|]���rR:� ��Ϣ�S�     ��0p��&�J P/l T%ǖ�6�8x<*� Tn8i���e�     ���)"��+�T�]�  ����d�)����X�>{9��      X�۟A�4� `�� �K㵍2�.���tP���Q�\�Kg      ,Lj}�ze9�J P/l �%�V2�����_�9>|pV:     `qr��g�+�V�[v� T� ���p��2FӶt     ���n�t �"� �d��q|1.�Td������      �Z�� ���; ��K' y��it}*�     �89E��� �
1p ��óQ�ɣ�gwx6�óQ�     ����t �b� �(��]q�M�r���t     �¥�� �"w �9{xj�<�>;�iۗ�      X��"�Y�
 `�� ����I�g]�`M=L���t     �¥v\: XA�  p��w�饔�ݻ��3      �"w��	 �
2p X��\_�����M��      ����~V� XA�  0�vq|�qz��;L���E�     ��Hݤt ��� 䳣��	���S���GΥK      �#�� ��3p X��qLf}�`�w�$&��t     �r�>"��+ �e� � 9G<8q��z�N��:,�     �4�s� �j�  ���t�¦m��?-�     �T�5p ���; ���>�F�3�����h�T:     `ir�"R[: Xa�  v��t������K�I     ���z; ��� ,��`��i�`�<L��ó�      K��q� `�� ,�+���̺>~��q�\�     `�r7��}� `�� ,���(FӮt�~��Q�Zo�     ���v �I� ,A��\q�����q6���      X��#w>' �:w �%yx2��K�3�B���q��]     �͔�ID�� ��� ��O9�]�� 
M�x��q�     �bR;.�  �	w �%�wt)����)��?9��w�     �P���g�+ �5a� �Dm��+�Q޽{�co�     ���v �i� ,ٝ���]q��p��Y<z<,�     PT6p ���; ���]��G�3�;<ŧ��Kg      ��YD�Kg  k�� ��;��C�.G�x��q�     ��r;)�  �w ��.ŽCWܡFӶ��||�K,      �#w� ��1p (���Et}*��QJ9~��QL[��     ��4"�L x:�  ��}�{���3�9z��q���3      VBjǥ �5d� P��Ë�u.=C޿�g��      �!���a  ��� ��)n?<+�<�O�����'2      ���� �U� ��d�I[:��ǃ�x�U      �R�y�- p5�  ������������'�3      VJ��/� �)w �pz9����ur1��۟EΥK      VKn}�	 \��; �������	�N�x��A�ɺ     �r��MJW  k�� `E�m�?�,���Yo�>��K�S      VN��J'  k�� `�|��,f]_:�
Ӷ���QLf]�     ��#��� ��3p X!m��g�3�/1����G1��     |��M#��^ ��1p X1Oqz9)����K��b8iK�      ��4s� xv�  +�{��s.�DD�r�u� c�v     �����~Z� ���; �
M۸spQ:6^���b4+�     ��R�z; 0�  +���M�������׷�l��     ��ˑ�Q� ��  +*���;)��O9��ȸ     �I�v�S� ��  +��r�Jg�F����� Ά��      O"�� ̑�; �����M����>�[��ܸ     ����E��� @E� V\�r���q��ެ���?<0n     x
y�z; 0_�  k�l8�;�3�Z���_t�c�E      �XΑ�I�
 �2�  k��g1���3�:�Y��� c     <��M"r*� T�� `M����O�#�\:�1����hj�     ��lX: ���; �����ó�P���4~����̺�)      k'w���s `�� �̝��8:�΀�vz9��nF�{d&     �U�� ,��; ���ݓ�:W��to�>�θ     �Jr�"�i(oZ{    IDAT� �R�  k��S���q�K��Z�t��=�      \]�y�4 �8�  k�|8���΀�q��Y��Ը     �Y�����  *f� ���^����ur��Ν����y�     ����qD�� @�vJ  �l�p�$n�؋���h���K�ۏ�l8-�     P�y�  �X.� ����|����$�_M�x�G��      s��iD�Kg  �3p ��p���?=.�+��ro���i[:     �i6,�  l w �J�\������3���'�����h=�      `nr�F$ǅ ���)  ���?��[7�⻯�*�E|��q�9�(�     P��z; �$�  �y��Iܼ�/?�t
,M�r���Q��K�      �'���i�
 `Cl�  `�r���'G1�x< �a8i����     ,HjG�Kg  �� �Bm����d֗N��:�Ǜ<���:      "�ȭCC ��� Tj����b��S�;�ۏ��S�     �j�v�} ,��; @�F�6~s�0��q�ԣO9~��Q|��qd��     X�i6, lw ��]�f�#[S�ᤍ7?؏óQ�     ���v�=1 X.w ���r���t<���a����1��S      6B�9: ,��; ��8:�;w�Kg�SK)���;w��O�D      ���D$�� ���)  ���#���G��N�'2����O�\m     X�4�N  6��  ���(~��a��6����0����q;     ���n�z; P��; �::��>92rg%�)����w���S�     ���f��	 �3p �PG�����G���;��b4�_��O�i
     PB�ۈ~V: �`�  ��b���0z#wV�������c4��K     �R�lX: �p�  ��ro~��Y_:�5�����g�}�     �����ݤt ��� ����7?؏���l���l�|�a���S      6^��� �g� @DDL�>���Gqz�"��v)޹s���(�>��      ��� +�� �?k�o�>�ǃ�)T��b�����?u     `U��0"r� ��)  �j�9��{'1m���Q:���]�>;5l     X59Enǥ+  "�� �����Y\�����;��ó9�ǻw?��      ���v `�X* ����o�?��-�j���9���>4n     XE9E��� �w  ��h��/�ۏ�'��)����a��w���t
      _!�F�Jg  ��N�   V_�9�p�$Ά����MӔNb���]�w�$N/'�S      �:9E��JW  |��;  O��� ��6~��W�ƞ%���s|��">}t)��9      �i6���Uc� �S9N�_�}?}����ϗ�aE���N��)      <��"�ƥ+  �?�  <�>����8���������]:�B�m���ÓA�      ���� ��2p ��N.���>����[/?W:�%J)ǽ�����yt�7>     �JN�g��  _�� �g��)޾s����w_�ݝ��I,���Q|��qLf]�      � M�Kg  |)w  �b�t�����_���|�`0n��'q6��N     �R���  �J�  �Mۧ����?��}��x��^�$�`�����Y<<Dv�     `���0\o V��;  sw1�ś���܊�}����jJ'q]���G�q��2��MN     ���z; �� X��#��|�����/?W:�'�R�{Gq��E�}*�     ���� \o V��;  5k�x��q�98��~��x�ś�������YL۾t
      s�S����  ��� X�����~r�x�Z����篗N�r����(>�?�Ѵ-�     ���0\o ց�;  Ku>�Ư?:�o]��y�x�ֵ�I+�O�.�     T.�.r�z; �� (�l0�_}�(^y�F��/��D)�|w.bf�     P=���ub� @Q'�8���7��{�=o��\4MS:�J���ώq��"�.��     `	>��>.� ��� X	��Y�{�$n���^}>���󱻳U:�
�q��.b�d)��     �I�tP: �� �Rfm�ŝ����K��w^�/޺V:k-�����E�^NJ�      P@�g�;� ��� ��ԧO��d��v�[/݌��|���#�יu}<<�gǗ1�v�s      ((�� �!�   V�d�ŝ���{x/޺�y�V������jJ�����q<8���q�\�     ��r7��g�3  ���;  k#�Ǘ�x|9���������x3^}�F\��.��t��Y<z<���aL۾t      +#�� �-w  �R�9N.�qr1���[7v��n�k߸/޺V�nq��6����a'm�      VP��#RW: �J� ��`��`�Ɲ����ݎ�n]���/ݺ���+��L·�8�����0c�v      �FΑf��  Wf� @ufm�Gq�x�[M��ܵ?�޿��^�lo��j�����q�\L��rm�J'     �&�l���  Wf� @������$_N"�<""�v�����x��nܺ��]߉[��bwg��������4����p�J;      W�S�٨t �31p `#��>N�>N/'_��ww��k����{��qmg;���_��?��lE�4O��ק�I�i�Y�I�i��Y�)��      *M��� �z3p ���v)κ��g��&���h�>��?�눈�s�)Gץ�R�l�     �"�>r;.] ��� ��RΑ�ї.     `ӥ�eD�� ����         \]���ݤt �\�        ��ϯ� ���        `M�n��Jg  ̍�;        ��J�A� ��2p        XC�G��t �\�        ���z; P%w        �5��Èܗ�  �;w        �u�S�٨t �B�        ��4DD*� ��         k"�.r;.� �0�         k"O�Kg  ,��;        ���,r7)� �P�         k M.K'  ,��;        ����8"��3  ��        `��H�A� ��0p        Xai6��}� ��0p        XU9E�KW  ,��;        ��J�AD��  Kc�        ��r�"���  Ke�        ���t�t �R�        ����"w��  Kg�        �b��t @�         +$���Ԗ�  (��        `e�HS����e�        �"�l���  ��        ���"O��+  �2p        Xi:��T: �(w        ��r�"���  ��        ����ȥ3  �3p        ((���ݤt �J0p        ((M.K'  �w        �Br;�Hm� ��a� ��a�β9� 
����$�2�}POR�' �*�l��{      (�ї��  �"p        (��KD��  �"p        x���k�
 ���        <Y_^"�W�  8�;        �e�#�k� �C�        <Q�}���� pHw        �'ɶF��z �a	�        ��� �_�        <An׈�U�  84�;        ��e��z ��	�        �/�٪g  ��        ���G���  � p        x���DD�� p
w        �ɾGn��  �!p        x�~�Y= �4�         �m�hK� �S�        <��{;  !p        ��ܮ}�� p:w        �����K� �S�        �Q_/٪g  ���        �^�G.��+  NK�        p'}y��^= ��         ��[�v�^ pjw        �;�˷���  �&p        ��l[�~�� pzw        �/z{o ��         _��-���3  � p        �����T�  ��        ��r�F��z �0�         ��}�� pOw        �O��kD��  C�        |T���R� `8w        ��˷��� pow        �ȾGn��  C�        |@�}��  0,�;        �;�F��z ���         ����  �$p        x��n}�� 04�;        ���v �'�        �A_/٪g  O�        �;���k�
 �)�        ~���٫g  LA�        �+�#�K�
 �i�        ~�//� �Y�         ?�}�ܮ�3  �"p        ��\^""�g  LE�        �ٶ��V= `:w        ���˷�	  S�        �K�KD[�g  LI�        �/}y��  0-�;        �_r�F��z ���         ��� �	�        "����l�3  �&p        Ȍ\_�W  LO�        L���٫g  LO�        �-{�z�^ @�       ����%"�� ��        �V�=r�V�  �/w        `Z��DDV�  �/w        `Jٶ��V= ��        S��K�  �C�        L'�і�  ���        ���v �c�        S�}�hk�  ~B�        L�{; �q	�       �i�~��[�  ~A�        L�{; ��	�       �)�v��{�  ~C�        L �� ���        ^�׈l�3  ��;        0����V�  ��        ���z�� pw        `\���� NC�        ���٫g  �Nw        `L�#�K�
  >@�        ���� �L�        �x�G���  |��        N_^�{; ���       ����yo 8#�;        0���DDV�  ��        �0��ۭz  �$p        ����v �3�        CȾG��� �L�        �߾UO  ���        ��e�"�R= �/�        ����  #�        ���޾V�  ��        ��yo ��        8-��  c�        �� `,w        ��r_�� F�        �R__�'  pgw        �t�� �I�        ���v �1	�       �S�� 0.�;        p*�� �%p        N#��{; ���        �i��{; ���        �)�D��z  $p        N����  x0�;        px��m�� ��	�       ����K�  �@�        Z6��  ��        ����  ��        ��m�� 0�;        pX�� �"p        ��}�� �	�       �C�� 0�;        p8�� �$p        '���	  �        ��m��o�3  ( p        �{; ���        �ad߽� LL�        ��v ��	�       �c�-r�� 03�;        p}}���� @!�;        P/{�v�^ @1�;        P�{;  w        �Z���{;  w        �X_/ѫg  p w        �Nf�v�^ �A�       �2}�D��v  ��       �"�zo �w        �Dn��l�3  8�;        P����  8�;        �t��"�^= ���        O� ���        O��ѷ�  ��        x���TO  ��        ��d�"�Z= ���        O��k�  L�        <Go���z  &p        ��{o ��        ��e�ܮ�+  88�;        �p}�DDV�  ���        �ceFn��  ���        x��]"�W�  ��        �e�� ���        ��-"[�  NB�        <L�� ��       ���}��[�  ND�        <D__�'  p2w        ���m�� ���       ����R= ��        ��=r�V�  ���        �]��Y= ��        w��� �4�;        p7��"�U�  ��        ����R= ��        w��ѷ�  ���        ���  |��        ���{D[�g  prw        ��r}��  � �        ��d��n�+  ��        ���^""�g  0 �;        ��]�G  0�;        �i�-٪g  0�;        �i}}��  �@�        ��d�"�V= ���       �O��R= ���       ����ߪW  0�;        �a}�DDV�  `0w        ��2r�V�  `@w        �Cr["�U�  `@w        �C��Z= �A	�       �w˶E��z  ��        ��z  �        �=r�U�  ``w        �]�v���� ���        ���z��  ���        ��Dd�� ���        �u��  <��        ���"�R� �	�       ���۵z  ��        ���ۥz  ��        �����z  ��        �Խ� �Dw        ৲�m�� �D�        �O�� ���        ?ʌ�n�+  ���        �A��3  ���        �A_/�  ���        �N�-�o�3  ���        �Nn��	  LJ�        �#3r�U�  `Rw        �o��"�W�  `Rw        �o}�VO  `bw         ""��m�� ���        @DD��v  �	�       ��H�;  ��        @�Dd�� ���        @t��  ��        f�[D[�W  ��        f� ���       ��R� �A�       `b��٪g  @D�       `j�]�'  ���        0���R�  �&p       �I�v����  �       ���v��   ��       ����}��  ��       ��r�UO  ��       `B�]�'  ��        0��׈l�3  �w        ���v  �J�        3Ɍܗ�  �Sw        �H��3  ��        0��]�'  �/	�       `�E��z  ���        &��[�  �-�;        L"�k�  �-�;        L ����  �[w        ���v  �@�        �}��   $p      ��*h    IDAT ���Fd��  $p       ���~��   �"p       ���� ���       ��r_#�W�  �w�       ��r�� �y�       `T���R�  �M�        �z��{�  x7�;        *�[�  ��;        �(�w  8�;        ��=�g  ���       `@}�UO  ��       �h�G��z  |��        ��Y=  >L�        ��۵z  |��        F�=�m�+  �S�        0�ܗ���  �)w        �[�  �$p       �Qd
� 85�;        �-n��  �iw        D��	  �%w        BF�k�  ��;         �%"z�  ��;        �-p �s�       ��� �!�       ��r�"�W�  �/�       ���~��   w!p       ���}��   w!p       �˶Fd��  w!p       ��� �H�        pbw  F"p       ���-���+  �n�        pR}�UO  ���       �I�VO  ���       �eF4�;  c�       �	e[""�g  �]	�       ��r_�'  ��	�       ��r_�'  ��	�       �d�m٪g  ��	�       �dr_�'  �C�       �d�  �J�        g�=�o�+  �!�        p"�� ��        ND� ���        p���#  �a�        p�����3  �a�        p�/�  ��        p���	  �Pw        8�̈�U�  ���       �	���g�  x(�;        �@�K�  x8�;        ��ۃ;  �M�        G�=���+  ���        pp�/�  �)�        pp���  �)�        pp�<� 0�;        X�-"{�  x
�;        X��z  <��        ,w�;  ��       �ae�w  &"p       ��ʶGDV�  ���       �A��v  &#p       ��j[�  x*�;        �w  f#p       �ʶEd��  O%p       �#j[�  x:�;        P��z  <��        (=� 0!�;        L�="[�  x:�;        ��v  &%p       ��ɶVO  �w        8���  �I�        G�="[�
  (!p       ��� ���        p ��  �K�        �m��   e�        p���  PF�        �m����  e�        pm�^   ��        p��  �M�        �� ���        � 3���+  ���         ��v  �       �d� ��        �@�  w        8�   p       �z�#�U�  �rw        (�  ��       ���  ��       �Z߫  �!�       ��w  x#p       �J�#�U�  �C�       @��{�  8�;        Tjw  �?�;        ��  ��       @!�;  �C�        ���  �O�        Uz��^�  C�        E�{o ��       @�;  |O�        U��  �M�        E<� ���   ���;�m]ɡ(Z�|���_���C'�-�,i-���`�     PbC�  _�       ��v�cl�g  @+w        ��a�  ��       @��.p ���        P��Q}  �#p       �� �'�;        T�,� �ww        ȶ�?  ���        �mw��  ���        �	� �!�;        $���T�   -	�        �w  xH�        ɶM�  ��        ����  �%�;        d��  �A�        ���G�	  Ж�        2	� �)�;        $���T�   m	�        �f�  ��       @��~�>  ��       @�M�  ��        ��Q}  �%p       �4�w  xA�        I���v  xE�        Y�� �Kw        �r� �+w        H�m�'  @kw        ȲYp �W�        ��.p �W�        �d�>�O  ���        ��.p �W�        �e�W_   �	�        �vcl�W  @kw        H�Yo �]w        � p �]w        � p �]w        Ȱm�  @{w        H�Yp �]w        � p �]w        � p �]w        Ȱm�  @{w        H�Yp �]w        �`�  v	�        �w  �%p       �� `��        2lw  �#p       ��mÂ;  ��       �Ѭ� �[�        p4�;  �E�        ۆ�  �!p       ��Yp ���       �pw  x��        ��o ���       �p
w  x��        'p �w�       �h��  �!p          ��;           -�       �h�V}  LA�          @w           Z�       ����U�   S�          Ђ�          ��           � p          ��;           -�          hA�          @w        8X��>  � p          ��;           -�          hA�        G���   � p          ��;           -�          hA�          @w           Z�          Ђ�          ��        p��>   � p       ���� �-w           Z�       ��L� �;�        p8�;  �C�          @w        8�w  x��        �p �w�          hA�          @w        8ZD�  0�;           -�          hA�        ��'  ��        p�� �;�           � p          ��;        .�  �)�       �h�v  x��        �p �w�        �T  ��5       @#�  �K�        )�  �G�          @w        �� `��        R� `��        2Xp �]w           Z�       @
�  �G�        	"�  �G�          @w        �`�  v	�        ��  ��          hA�        B�  {��          hA�        "�/  ���        � ��  ��        �w  �%p       �w  �%p       �w  �#p       �� `��        R� `��        2Xp �]w        H� `��        2Xp �]w        H!p �=w        �`�  v	�        ��  ^�       @+�  ��        �� ��;        d	�  ���        Y;  �"p       �4w  xE�        I;  �$p       �,w  xI�        i�  ���        ��\  ^�c       �,a�  ^�       @���  /�1       @�  ���        ���  ^�       @�;  �$p       �4w  xE�        Y,� �Kw        H!� �W��        �w  xE�        Y"��  ��       @�� �3w        H%p �g�        �)$;  ���2        d� �S~�        �("�O  ���        �ɂ;  <�        �,� �Sw        �d�  ��[       �D!p ����        UT   m	�        �w  x�o        2�w  xF�        ��  ��        EHv  ��e        �d�  ��       @���  ��       @���  �#~�        �M�  �)       @���  �%�;        $�  �2        d� �C~�        �M�  �)       @���  �%�;        $�  �2        d� �C~�        �M�  �)       @���  �%�;        $�  �2        d�e�a�  ��       @�� �ww        ��  ��/        *� ��d        (w  ��/        *� ��d        � p ���       �@� ��d        � p ���       ��"� ����       ��w  ��/        
��  ~�K       �
��1��
  hE�        U�� �~�        PE�  _�!       @�;  |�        EB�  _�!       @�E�  ��        �Xp �/��       �H� �?d        �"p �/��       ���  ��C       �"���'  @+w        �Q}  �"p       �21FXq ���        P)$<  ��1        T� ����       �P,k�	  І�        *Yp ��       @�� ����       ��"� ����       �R��  @w        (!� ����       ��"� ����       �T�a�  �w        �k�  Ђ�        �Yp �1��        ��"� �1�        P/��  ��;        �E�  c�       �^�x  `�;        �� �C�        �bY�O  ��        P-�1FT_  ��        Ёw  �       @!�  �b        h ;  �       ��E�  w        h B�  ~�        Ёw  �       @� @�        �w  �       @��1��
  (%p       �.B� ���       @�Z}  ��       @!p ���        �E� �6�;        4a� ���       @� �8�;        t��y  �6?b        h"�  \��        ڈ1B� �u	�       �+�  \��        	�  \��        :�� ��	�       ��� paw        �$$=  \��0        tb� ��       @#w  �K�        �D��  ��O        ��� �E	�       ��Xn�'  @	�;        t�Xp ���        �L� �(�;        tw  �I�        �Xp ��        �Ͳ�1��
  H'p       ��B� ���       @G˭�  H'p       ��bY�O  �tw        �H� �	�       �!�  \��        :
�;  �#p       ��b�U�   ��        �Q�!� �Z��       ��X�/  �Tw        h*�[�	  �J�        ]-� ��;        4e� ���       @W� ��;        4w  .F�        ]���  �"�~       ���� �u�       ��Xn�'  @�;        t�Xp �:�        Иw  �D�        �Yp �B�        Иw  �D�        �E�2  ���        ��� �E�       ��X��   ��        ��� �E�       �9�  \��        ��� �E�       �����>  'p       ��b�e�>  'p       �	�r�>  'p       �Xp ��        0�  \��        f p ��        0�X��  �pw        �A,�  N̏        f�ܪ/  �C	�       `!p ���        0�e��   %p       �IXp ���        0	�;  g'p       �Y,��  pf~�        0�e��   #p       ���z�>  #p       ��,w  �K�        	�;  '&p       ��� 83�;        �dY�� ����       ��,k�  p�;        L&�[�	  p�;        �f� pNw        �L,�O  �C�       `2���'  �!�        0�e�  ��/        f�ު/  �_'p       �	�"p �|�        0�e��   ~��        &��  ��	�       `B�ܪO  �_'p       ��2F��W  ���       ���� p2w        �T��O  �_%p       �I�w  NF�        �Z�  ���        &�:ƈ�3  ���       `Z1�b� ���       ��b� pw        ��w  ND�        ��O�	  �k�        0�X-� pw        �Y,�  N��        f����   ~��        &�� �s�       ��b�U�   �B�        �[�  ���        &���. `~~�        pV� 8�;        ���;  �M�        '��  ��&p       �3�� �	�       �b��1��  ���       �;  ��    ����Ǯ��������)�EY6eS�eE�D�X��4
6.p�"�Vۥ��v*��VR��O��-�,���z-k%Q�1��P$[�g�9�{^�V?�H�{9��\   ��w  X.�;        4"��z  <�;        ��w  N�        �p� ���      ��Ml    IDAT @+2#:W� X.�;        4�w  �L�        -�]p `��        А�]p `��        А��  ,��        Z�!r `��        И��	  p*w        hL�� �B	�       �5�� �e�       @c�""�g  ��	�       �9��#  ���        Р���	  pbw        h�� �%�       @���z  ���        ��Y=  ND�        Mʈ~�  '"p       �Fe7TO  ��       @���TO  ��       @���'  ���       �U]�}�
  86�;        4�w  �D�        -� � w        hXvw  �C�        K� X�;        �,3�w  B�        ��~��   �"p       ��e���   �"p       ���c�  8�;        4.�!�B  ,�W�        ��P�   �J�        +���z  <��        V ��z  <��        V@� ��       `���D�  ̛�        V�w  �N�        +!p `��        �w  fN�        +����!  �˫U        X��7�  ��        �&�X�   K�        +�;  s&p       ��~����  �$p       �UɈ~�  �$p       ��I�;  3%p       ���~S=  I�        +�;  s%p       ���.�� 0?w        X!W� �#�;        �P���	  �w        X��  ̏�        �(���W  �7�       `�\q `n�        �R�� ��;        ��� ���       �Zu}D��+  �kw        X1W� ��;        �X�c�  ���        �lp� ���       ��e7Dd_=  "B�        ���X=  "B�        ��öz  D��        p� ���       ��e7Dd_=  �        @D���	   p        "r� PO�        �� �,�       ����Ⱦz  +'p        """W� �%p        """{�;  ��        @D� �'p        ����W�  `��        ��r�VO  `��        �ײ�TO  `��        ��r� PG�        �^v�X� ���        ���;  U�        �7d���  �J	�       �o�a���� �
	�       �oɈ~� �
	�       ���a[= ��        ߑ��z  +$p        �#�1"�E  \,�@       �Gr� ��&p        )�m�  VF�        <��  \4�;        �h]�}�
  VD�        <V��	  ���        x,�;  I�        <V�����  ���        x�̈~S� ���        O��� ��!p        �(�m�  VB�        <QvCD��3  X�;        �T�� p�        �S尩�  �
�       ���~Y= ��	�       ��ˌ���  4N�        K��	  4N�        K���	  4N�        K�cD��3  h��        8�\q ���       �c�a[= ��	�       �c�~Y= �F	�       ��ˌ�7�+  h��        8��  ��;        p"ݰW= �F	�       �����n�^ @��        ��尭�  @��        ��	� 8w        �Ĳ#R~ ���
����       �!#�M�@+@c� 4%#��       k�öz)p�)w �2M�m       E�s��J �6 ڒ�m       &��~S�V�w �"�1�g      �r��i% h� m�:�6      �$p�Z��1l 4eJ�      .RvCD7Vπ��t� �Ń��t�m       �w(��� �,� h��Wo       X�;ԙb��)l ���n      \��ǈt��h% h� mI�6      �
��C� h� ��l      (��^�X��.�7 �YД�&�6      �9�!G�Z	 ��@S��<�       Jd䰩듓� 4E@[�i��       �V9�UO���B+@S� �%c[=      `�����4\�̱z �%�; ��      T�.��T�����x�CW�h������      �BݸW=V�ͧ��; ��      �Pۈ���*w�P/@3� ��w      �J�E�c�
X�m�� �w Z��       źa�z�ʃ]�K@3� 4dʈp       �X�Z[�HC�q��f�h�[��cDd�      ���.����E9�����f�hƯ���7k       3����E針�p 4C�@3��]�      ��nث� ��;4 4C�@3�m'�F      ��������
]i& h���f���       s��+�p:� �Ќ�G.�      �I~�a�e�w ��1�Wo       ���"��z��A�  8+w ���]��       �7�W=��;�; ��Ў�	�      f��p�v�� �w ڱs�      `v�>��W@�v]�; ��Ў��       3��+�p�r7	�h���f�ެ      �P7��\e�WO ��"p�.�      �S�G���ЬGh������      `�\q�s�[�h���v��      0[9
�Ἰ�@K� �ç�      �+��~S��4E�Wo ��"p��L�      f�\q��0M��� 4C�@;��      �X�{��3�Ew �!p�%w      �9�.��T���dN�� ��hF
�      f���'@�:�h�������       <Y{��3�)S�a� 8+w 2=W�       ��Ȍ��+�)��]��  gE�@K�       ��^�hKƥ��W# ��; -�R=       ���a��%8C��_��a� 8^%Є[��W���      �qd���;���W�Vo �� p�	��x�z       Ǘ�����=�V� ΂��&L)p      X��7�WπfS�� �	w �0��I      X���'@3�~�� �	w �0M�M      ���W=�1ew�z ��; M�B�      �4��X=���j' h���&tޤ      ,�+�p6�]\��  gA�@��w      �%����	І����; ��	�      �(��~[��o
� M�Ј��       ��+��즌�� �,�h��      `�r�~y�8�)���  g��B ����^�      ����a�z,ZNӵ� p� ��w      �E�Q��$��� �,�h��       K��&"���\S
�h���F��      �t9�WO�Ś2� 4A�����˥��       �	���2�͍�?<�� �J����_\q�      �]�o�W�bݿ�ߨ�  �J�����\��       ��p�No�$p`�� ,^�\p      hD{!k��麝����J���<r�      ����z,Үs$����x����      �!9TO�E�v;GX<�; ��w      ��d?Ftc�X�k� �Y	�h���       8[9�UO����X<�; ؽ\�       ��Ս���3`Yv�#� ,������	       ���"�m�
X��� �Y	�X�.nVO       ���xP=�e�]��  �J���M�;      @�r�Dd_=�w �O���]�����w       p>rܯ� ˑ�SV� �g!p`�r|p�z       ���I�7?��׫G ����l�N�      в����+`1v��[� �Y�X�)�       ��6���q=|8h) X4�; K�M      @�r�Fd_=!� ,����˗�       p�2rt��c7MZ
 M���yS      �
���%�x�z <�; K'p      X�����W��ej) X6�; ����To       �b�+��T��; �&p`��W/       �b䰍Ⱦz��4ݬ�  �B��b���݋��w       pqrsP=f-C���	�X��>��{��;       �8ݸ~TO��B���P= NK��b�}���       \��"�m�
�����U= NK��b�v��      `�r<�� �6<��Wo ����XSī�       �x9l"��z��ԇ�� ,����ʈW�7       P�s�kw �K��rM��      �J���'x�)oUO ���
���x�z       E2��܁��I��b	�X��w      ��ƃ�	0K��^��  �%p`��|��6"nT�       �P�G{�+`v2��� �� ,�?歈��       �JW�Ủ��Xw )��]�      �z9l"��z�Kƕ�����3 �4� ,�Qt�Uo       `��+��mG�� ,������	       ""r܋H)��.�� �4��`�2�v�       �"#GW��M�
 J��R��      �׺q?"�z�G���' �i�X���       ������+`6r�� ,���Ź��Gۈx�z       󒛃�	0��j� 8�; �����      ��d�����0SN�To ���8]���	       �T�;DDDF܌���O| �8w �{�z       ��^D��3`��n��j� 8)�; ����]�      ����q�z��Ç�~X� NJ����"]p      ౺�ADd�(�������89�7_       <^v��^�
(7��� pRw '#^��       ����z���� pRw �ֿ���)�Z�       �-�1��g@�I��	�X����7�7       ���R��5�nWO ����(�._��       �2��}�(�7�|�Ѷz ����eI�;       ��;+��c��U� ����(ݴ�      pl9�G�L���ؾQ� N�+7 e�\p      �2#ǃ�Pf�t��E��,w�'       �,�� �R�U�$p`Q�j`1��ٯ^����;       X��"ǽ�Pb��� pw #��Wo       `��ͥ���p�r��7 �I�X�.�7�7       �P]9���M߯^  '!p`9��S=      �����	p�2^����J� 8.�; �1E�Y�      ���n���3��僣7�7 �q	�X��V       `ٺ�+��Q?��z ���E�����U�       `�r�Dtc��P9�~R� �K��"|~���W�       `�\qg}��� p\w !NoVo       �9n#ҍ5�#c�S� �K��"Lw       �HFn�G���"o���; �8� ,BF��z       ��ƃ��O����A��z �Wh ,�.�      p�2#GW�Y�i�{�z ������+�^��      @[��ADd��(?�  �!p`���x�G���      @c����W������ �8� �^��f�       ��m.UO�1M��� �8� �^F��z       ����a�z����a� 8�; �7e�U�      �v�+���ҵ�W�U� ���0S�]=      �ve?F���p�2�}G�=�; �v烏��O�w       жn{X=���92��	�����oF�X�      ��}y�}S=�U��� ̞��Y�.��z       ���;����O�7 ������Wc      p1�߸�N���� �i� ���;       �۸�N�2�����+�; �I� �[
�      �89��N˦n�oW� �'�0[7�э��Y�      �u�6��'�9z��  �&p`��ީ�       ��䰍���p.��V� �D��lMS��0       %��+�4j��TO �'�0_]�]=      �u�a�w�4���� �$w �k7�S=      ���6��Ӟ��u���V� ���0Kw>�hoU�       `�r܋��p�r�?rt���0K?�y;"6�;       X7W�i�.�Wo ���0K�����       ��+�4'��w fK��,M9	�      �W�i��v� x�; �4E
�      ���"���gg�~�~�Y�`~��WcF��0       3��m�G���8��o�N� x�; �s�ߊ���       �W�iδ��� �Q� �Ov�VO       �o��6��G���M�;� �Q� �N�$p      `vr��;��Q� x�; 3$p      `�2rsP=�H�U�  E��������       �R7D���˜^������� �m^i0+/u�y3".U�       �Gʌ���6M�q;�[= �M����v�UO       �'�6�Wπg6u��z |�P=  ��.�_e�fo;�q�7����f�c3�1�]�]F�_�	:���h7��n���ރ�q��Q|�Ńxp�+�       ˖�mc��慎�3�I�������|/b����}W6q�`�����	��w1�}l#"�_��{���/��>��~q?&�      ��q/�ާ�Q�8�)�w�7 ��9��l���=�̏#���]f\���.�ǥ�1�^�<<��ǟ݋�|�E|q����"      @��w]qg鎆�ϟ�����g�C �+.�0}���n7��Wn����A\;��R���.�_ُ�W��ӻ�>����޹��      ���q����cZ,V��ßE��� _�0G��=_-�^_��/\ދ����p�?���w�?������c�;      ���0vw?���v���C�����������}/^=��W�#g�3�^�׿x��7���{�-       ���^D7F�TO���x�z �!�; 3�?�^�źvy/n=)�����H���x�ֵ��O�Ư�Y��I      �}y����3�Tr�ީ�  h&wRX���������;�{�!^�q9������������I|z��      ໎>�ǈ���3�4���ϟ�����g�C  "b��RX�a߫���ˌx��A��ʵE������|5n�p�#�      ��t���	pZ�.V= �"p`.~^=��5]ܹu5^~�Ң���ǝ[Wc��      ~/�MD����r��6 �e 31�I��ϕ�����>VO9�1�x�Z���      �F��\=N'���	 ��; ��|��6"|�U�^~�R�v���^v}?�y5���W=      �������Y���w�7 �W�*� X�O.���7�ˌ�/����    IDAT]��TO97��޸/?�z
      0���Ch�޸�'���{��5�����u��޽}������1v������461c443ʌG�0�W#ED��`��H�m����m"�r��͈DJ�&b2�}�Z�V�����E�>�aw�CU=���Hv�v��W�vתU���� ,w @�X�NW����_���S�ų7�+ۑR�      �6W�YJ)�e��S�3  ������WȰߍ|���wk���+��=���      �۵ౕ��ӵ  ����J�� ���A/~�����K��[#w       RӍ�ݨ��%E�p� �0p���_��("������n��^���z����5��^5r     �u�[��,�Rʇj7 @��; �u���j7��v7���.D�xs&"��A�te�v      PQj��z���<R������� � ԕ���������>�b��]����l��       *j����\:��3� ����J����������u��!�{f3.�kg       �4W�Y*%�Gj7 ��; ռ���\����������{����F�v      PI3�3-�E)�'j7 �WN T3o��"<�m)������EJ���nz��)      @���߬]�$E�h�|�[���f�@5%��x|�n�����v��xT�&����      �����"��X,������� `�Y�PM*�˦Ӥ���/D��%���;�ޫ;�3      �R:��(��� �7�4 ������b����<��^݉��'�=�[��za�v      PA�o���RhJ��� �7w �z�߹/�/oǅ�A팥�¥���jg       �.E3��g_N�õ Xo� TQJ��xt]?5)E|�s���x      �&����X,��K������ `}YVPG)/�N��z�x�UWNS��ċ��kg       ���2h:���� ��2p��=s�;"ŏ����5)��>��&�NY9�l��֠v      p�R���B[.�3� X_� ��~���N���KW�c�߭���^�����c      �n��'>��J���	 �/�* �]i��xw�w7��ΰv�J�v�x�7�      `ݤN/Rw�v<TJ�W>�͝� �'w �_I/�N����x��V팵pqk�<~      ����T;�^�n�~�v ����s�̵�\�(�y��Ӥx�s��4�H9//^ގ&��      �JӉ�sŝŕ">^���d����G�������^����?E��m�y�     `�_q7�ba}�v  �ɫ# �W�O�N��v7�qygX;c-]�݈a�[;      8O��4p���Oĵk.�p 8W9��vo�Ӥx��N팵�R�K�������j�   �NJ>�m9�M��"JDD��˓z�Ž��;K���a|�?x�_o�����SDJ��ٻ�����1   N�ߌv:�(m�x��s�����[���b����|��/�(����{��v���R��F/.l���v
  �
*�������˽?%Gyӯ���C�gX|ʚ�C�tw�D�;�O�� ��?����E���  �4�hۑ'�k��[���υ�; ����s�D��ka�iw��v��3��.mŝ���C�   <T���������w�~o��hW�W[����*��}��ߖ���?�0|词�  �I�mDL�yV;ޠI�g#��jw �^�87)�_���[u�ﹲS;��^'.�n�����)   �<0\�m��F����s����������:�O�����9�u��:��1|��b<  ��i�;��7jg��R>QRDr��sc��9))����+;�뺢�H���7_�D��?   ������<^�w}�}���Si���}�O�[��m"��������t\�  VV��#u�Q��)pOJq��+���^�7��n`}�p.�{��~��x�vo��ыg��3x�n��+6�?��N  x'����x�>�7jwy�ww�J��!�[G��d��=�7wG���  �PlG��;<�ݼ�OD�p~�8'��x��"^��];���za3��Lb�~   ��ܿ�o��윏r��Z۾�>=p���|:�-  ��JM7Ro#��1,G��g"��jw �>�89�/�T��]�݈�����Ӥ�za#��Q�  `������!�Kr,��O�����0���{��1��;  P_3؎v6	OAcQ��()"yC�saj��{�z��g�ݏ���)�v������K�E�s���7\q  �^)'����e�y�v�;k���{7R�d����   �)OGQ�^���4i������jw ��m��]�z�#aܾP^��eܾ�&���a���?  ����;d���}Cv��D���\~O���7���vN����  �hz��NǾgga�����0p�\�p�Rz�v�m�qigX;�Gtew#�nF�=�  xL%_co�Ǻ�����x|��CN~u"E�&R�w����<  ��H)��N�ɭ�%%��F�S����V �\*�CV��=W�k'���&.��ۇ�S  �E��7��K;s��E�(m�y{�W'����7�߽I  <��F���v
D��hDI�� ΜwR8SW�}����߆�9���0�{u�v�i:�����(�&   "�/���(�ɐ=�"J�]��to螚�� ���m  <\ig����3 ""�4�������w�; X}.�p�>���I)�{f�vO��m��� n�N  �[�Q��ɐ�evXn%"ώ��<��y`���Gj�F�  �=�Ӌ�݈2��g꛷�OG��; g���3դx����pyw�nS;�'t�¦�;  ����'��{�فՖ���ߟG�{��=p����ݐ  ���w�=8�Op�����"⿮����n( g��_w�M{ߍ�K�S�]�R|�{.E�c������q  �����v�������N��w�яH�� �u���Ljg�������K�^��.`�����y6�$���Ջ��+��;  ,���٧'���xT%�����:�:w/��]y ������F��v
k-�\�h?���.`��pfJ�WRy�g�Ӥ���Q;�Spqk�ib޺�  ˠ��7�� 8M��2o#擓���W����wW� `u��`;��v��\��Sa��3p��4�|ƾ���6]o_)E<�=��n�N  ޢDi��>�(>�
��������ԉ���Gө�  <��ۈ��#��>SO)�r� V�gUp&����Ws��aY]Q����}��4�䯊ɴ�����Q;  ���F�O#�YD�.u"u�'�� `�vy�_;�5VJ�E�u�ƿ�Wwj� ��\p�L��J��ڞ��iܾb��Nlo����U  8w�=���,��F�F��<.u���w�  �$�_���'�SXS)�^�g~."���- �.w �Fi>QjW��n���;������Cw  8%�#ڙA;��Je���4�{��S��ܯ  �E�v�����SMI�w ΐ�; ��G��u����t�uwyw���+��� �v� r�  ���O.�_i���.8_y%ϣ��ǿnzo���  ��D�oE��.am��k �ڜ� �Խּ�rD���Xg)E\�٨���4)v7��3  `%�v�� ��h�����Ӹ "Ϣ�ƑoF{��h�7"OGQZO� �ښ�VD���`m������׮ `u����K�sW��K;����*{fg�FG�3  `����J�Q�vQr�"�%Q"����C#"R�ӿݽ1� �s�R4Ýȇ�j���J�s�LD�O�K XM� ��R�/�nXwWv]o_u;��v����8  �nJ;;�Ϗ"��� ���(�I����שs<v�#u{��� �:H�aD��Nk���R*�w Έ�; ��k��?+�W�c�]�İ�b֪K)bw�7^��N ��S��+��#W��Ci���Qf�h"u]w ���w#��#�s�9_%�/D������kj �bR�s��������[��	  �0J;�<E;���w#ފ2;4n����{�܎v�Z����GQZO�  �Ӗ�n���SC�z��� �&�8U%�����A7��������~t�m��x  �Q��Σ�O����� x�<�2�E�D����{w�ۏ�T�  �^3؎v>�A�]��~)"�m� V�� �����g#�õ;�����8G)E�� �:)\~�����(��q;�2)9��0���㿗{�  <��D�߮]�z�D�  V��; �&���זj��&.;����~�  8[�=Bފ���!dB,�>�t��h�7�L���  �R3��o�[��g>��/Ԯ `�tk �:R�_�H�z��D�?�����GJ��. ��S�<�le~�g�s 8/�4r;�8���"�����H�g ��h�;��7jg�FRJ�No���k� �Z\��T����lF�O��Xg�v6j'PA�I�5t� ��W�<��A���ȣ�(��v�u�gQ�^�<�;~���N��4"|�  &u���~n������ ��q��S1ߜ&Jڪݱ�����;�3�dws��?  ,��΢�'Qf�����`Q�6�le6�H����a�n�v  ,�f���("r��D)铵 X=.�p:J�B�uvigX;��v6�0 ��Q�i�ɝ�k���(ӑq; ��d�oܿ����?  ��t"ܦ���T�s����Gjw �Z\p��}�;�t��E��Ӥ��5��AE�~'z�&f�+  ,��N��&Q�G�� ��7_v��/�wz��  ������0"�k��&J�."�}� V�� <�go�/���XW���4�v�mm��-  ���y䣃�K�7�Ǉ�� ���F��"��]v �H�vkG�FRI��n `��p
�j��K;��	,��~�  �?j�E�E��p�N.���~����GQ\� `ͤn?R�ϒ9'M|����/�� `u��t�_o"�/��XW�nl��3X �C� ��mG�F� ,�<�2=�<�;�OG%׮ �s�v�<��"�ݍ���; X^� �T������jw���[��	,�A����v  ���#OG�CA�v �E�E9z=ڃ�F;�evh� �jk:�[�+X95� �+( �Jj�j7���<`�w  �T�2�D>���kQ�^�ȳ�Q �d�i���h^�|x+�|�v  �����x*8g/����8�� �>_;`]m�1�ujg�@6�  ��2? �n �*z����N���  X%)��n��AJW��L|�v ���� xbW�}�Ǣ����XW]o�M\p ഔvevx<f/�v ������Qf㈦Mo#Ro�܋ `��n?Rwxr� �N��+��� `�yG�'֤����w�d�ߍ&��  ,���L�ю�#����}�� ��<�|t����'�  ���n��q�R�O�n `5x��+)~�vú�tc����`��t��  <�e~������ND�Վ�R��''_+�"O�D���Q  ��Ri�U��U��/~���jg ���x"W^���%~�vǺ��z;a� ��(�,���Uڛ����(m��8�h/��(�CO; `�4�͈��9S���/׎ `���D:���nXg�y�a�R  <Dɑ��hG{���Qfc�< xR�4���ɇ�nGi���  ��h���#Xq%���n `���DJI�V�a]���:�3XP�  �I�O#ފ��(G�G�y�$ X!%��0����Ȧ#  `��N?Ro�v+,E|��Ǿ�S���f��c�������jg�W;����FJ�+  �.����^�|x#�|�v ��<�r�����[Q殺 ����ND2㌤ƅ�/�� `�y��ckr�V�a��l�k'��R��\q XO%�|��f���k� k��kr><��^���f  ,����᬴�_�� �r3p�	�/�.XWMJ�5p��w6�uj'  p�J�G�ܹw-6ڣ�I �]y������N�<�]  �z��8��OǇ�n� �3p�<��~2"~�vǺ���iR�ܠo� ���(���ȣ�(�qDɵ� ���Qf�ȣ�hG�Qf��;  u5�݈��gN_��x�ʳ�P���e��cɑ��nXg;�>Aϻ���  8+%G��N���t� �Q�E��v� ��RӍ�߬���J�/�N `y��J��mox��n�s� `Ք�4��h�������N �Vy���f��� p���vD��E��gk ���xdW����"�}�;�U���F�en���� `5�e:>��~#�|R� 8+�Q�Û�_�����k �.R�f�S���Ry��O_�p� ���; �,5�˵���f�vK�iRt;^� ,���"O�D{���k� �NJ������;��   �^�#u��3XA%ů�n `9Y>�h^�ލ_���ζ���	,�^��< ��RJ��a������(�qD��
 �+G������V���v  +��)�-E��� XN^� �H�\}���l�u�9��N`�����	  <���'��_�<��g�� �S�ȇ7�߈2�DD�� �*j:�[�+X5)����W�v ����G�4����Ӥ��yt}� X�2�D;�y��Z; �h�i�ɭh�"OG��  NW�ߌh<Y�ӕ�ޫ� X>�O ��?���(�˵;��Ơ)ծ`��\p X<�D���Gi�[�v ��J�����w��y�"  VF�f�[;��">_���c���j���#b�v�:���<����2 `Q�<�<���k���D��v �r��8�h/���(��A  ����E�m��`�4��~����� `�X>��R|�vº�tk'�dz�  Օ�4��ȣ�(�qD��I ��j�"ތv�e6�] ��k;��95�i�# X.�O ���\�.��O��Xw.��:�T; `M�(��hG��oD�� �(�"OnE{�Z��8"J�"  �QJ�wkW�B�H��� �r1p�Mc�jD�kw��^��^חl��  ����Q�{�'�#�v ��J����k����b� ��I�A��v�"�O<���S;��a��;K��j'��-��y�N�w �3W�<����ԣ�#J[;	 ��F�D{����=�. `�4�݈d^�i(Mt�֮ `yx�C]��_�`D�H�u7�wk'��w �3S��ȇ�"������** �����}/��ND��<  Aj��o׮`E�h�P���a���u�W#�B�����;O�i�� �T�ev�h/��(�I�" �ǔ���ǯg&���y�   \�oFt��3X)Ň/���T���`��C��J�r�
\p��u/�  NEɑ�^���ȓ��` ��;��^�E>���� `�5��p�S�)�ޫ�# XVO ����/_���ݱ&�]_�y2M�& ��(yyr;ڃעLG�k' ��2�D�G;����� `����U;�U���k' �,� x[9�Wk71�wj'��:��; ��(�,��ȣ�(�È(��  �^{y|#��Cw  ޢlE4�>��I)>z������3p�-���?ۊ�_��A�F�<9� Ͻa�x?�|R; ��vj� ��H�/Ԏ`�uJ��v �����(��_����D�y
�� ����Q����  2t �MR���Y;�%�D��j7 ���x;_��1w��y; �;)Qf�ю�"ތ0� x{��  <��D�N��Y*?y���3 Xl� ���k�~)Ry�v)El��4,� ު�(�q�{�'�#�v �r�7t���ծ ����^�]�rKm���� ,6w ޠ��W#�ǭ��׍d��SH� ����Gю^�|t'����  �S{y�o� ��R���Q;�eV�k' ���x@I%�wjWplc�z;O��R; ���F�܉�`/�� ���E  ��� `�5Ý�dzƓI)~��O��kw ���� �.��]    IDAT���>�������;Oɾ Xc%Ϗ��(�qD� ����{>�e� �NR�`�vK�i�_�� ��2p������nྭ��;OǾ XG%�#ފ|o��U �y(�����vDnk�  pRo�;������� ,.w ""�k߹�Z��c)E{�<�R�� ��q|����}>�� ����0��^�ɝ��):  ���F$4�@���?�P� �W DDD/�#b�v��n4M�����o �Aig\l?�� @DD�(�q�{���Q ��R�`�vK*w���n `1�)�߭��}��yz%�� X]%Ϗ���}� V�2=�v�Z��(��U  +)�6":��,�r-�# o� ����GK��>-����;O�a, `��b�a; �r(9�����E�y ����N���R�K�?=��� ,�* ���?���m�yz� �*q� `�6��V�#��  VMj��[�3XF����	 ,w�5��W�|PJ���ܗRİg���+� ��{�v� VG>~*O;���ծ ��4���N�v��W����d�v ���`ͽ���Ո�R����n4M��  U� ���(�x?��(y^� �S�^�4K�����jg �X�� Xs����n��6��s:rv� X>��� ��2�D�G�܉(�v  O��Dlծ`����f� ��;��r�/(��x��h���Sb� ,�{�����  k�D����E��"�{[  ˪�oEt��3X*���}����+ X� k�I��""����6��	���� X���.� Qr��ף��# �2�/�i�*�ԛu�/�� `qx����ʟ"�Wjw�FMJ��w���WJD.� ��m���v  ���!��(y^� ���t"�jW�DR�ߨ� ��0pXSwv��"�j��hs؍�>��͹v ��+9��A���(�q�  ];�<ڋ<�Q�� �L��VD�_;����+���Վ `1���߫�[mz�X��v `����E�D�,  <�2;�v�y:
�% �G3܍W�x$���# X� k�W�����X��jsЭ���p� X�D���/�O"��  �P�Q�^�v�e>�] �#HM7�`�vK���R�u�F ��Q.���H/$�9-�	w ��r��f9z=�� pJ�<��h�7��y�  �E�ߊ��kg�R��.z��; ���`ͼ���_���[�{��u}i�t�� @Eev��^������ `U��ȣ�ȓ;>P	 ����n��ǣI�S� ���� ��Q^-����6��	��\���W�Gю�� 8We6>~r�t\; ��HM7��N��AJ�|�c����3pX7)�~����W;��; p�J;�v|#��͈<�� �:*9�ѝhG�QZ�I Q�oFt�3Xt)�۝��kg P��;�y�7��R�O����m]p����G2 g��y��[����v  D�Y��ݧ
y� `�t6.D$�5�Y��[� �˫�5RJ����&������� g�ް}�e>��  oQf�ю���k�  ��D3ة]��K)}��g��C�; ���`M<�ϯF�k�;x{[�^�T��U2�� g���G�G���  ,��#OnG;ڏ��j�  p"�6"u��3Xl���ߩ@=� k�D���;��5t���5�� �i*�/`N"�� �G�g����'�#���  A3܍H�k<\I�7#���`M� ���u�4������9m3��SRf�h���  Xz�>�9;�� @j�G��)��\ze��� �a���M����[����R��[;��fWU��S�Y���'�"J[;  NGɑ'���Gig�k  �Z�#u7jg������� �a��J�o�n��6�h�T;�RJļu] x2%�#ފ<ޏh��s  �l�Y��' T�w"R�v�D������� �?w��«��@�x�v�5��N`�� O��ȓ;�G�Q��5  p.��������  u�&���,�T����Wkg p��V\[�?�����;�mf� <�e:�v�e6��R;  �Wi��btx+"��k  �N��#�6kg��R�|�v ���`�]��?ߍ(_���;3p紹� <�2�D{���ND� ��V��k��q� ���v"R�v�郗>�?];��e��º���#b�v�1�F�q`��e� ���΢߈<�Q\� ��r�;юoD���1  �#�h6.֮`A����n �|���k݉H�_;�w�z;ga67p �^��ȇ�"��#�i�  X\�4�h?��AD��5  k!uz��۵3XD)�x�c�ܩ���1pXQϦ��G�������l�k'���殰 oRr䣃ȣ�(�I�  X%�� ��~ 8�`+����Y�iw�_�]��1pXU����	���\p�l�����a���(S�' ���y��ȓ��� �V���B���fMi�V���� �
���_��H�3�;xg��^t�T;�4��! Q�Y�F8  pj�?<�H  g��D3ܩ]��I�᫟������0pXAMi\o_���s�Jq� �^n#ގ<ޏh��k  `��6��ȇ�|� ���F��v&���k7 p>�V�s_����j����F�v+h��(�v PG�|tprQ�v  ��2�D;ڋ2�� �4�݈d��}%�K/~��f� ΞW  +���DĠv�Ӥ�����s� �S�E{�ez�H ��(9��v�㛮� ���D3�X���".N��Wjw p��V����?#������m{�R�
V�t�i �NJ�G;���fD�A7  ��=r� ���n?R��n�K9�^���g��BG�������mo�k'���3�6 X%G�܉<ڏh�j�   '����-�� NY3؉h��3XM�ЕO��O�� �l����כ������lo�j'���sw Xuevxrr�v  ��2��� p�R�fx!"<&�c��|�v g��`E<�7W?�">P��w��4����r��l�: ���N��G��v  �k�  �.uz��[�3X�.�|�b� Ύ�;��(�Ok'�h�\o�Mf��	 �i�m��[��7"�v  ������G�Oj�  ��f�����`���گ�� ��������?�~�v�fwsP;��sq� VJ�2�  �2+'Xu� ���/D$�7"R��k7 pv|�XM4߬���I)b�w��d��N  NIi�юnD>�F0  ��\s 8%M'��n�
A�>p���� �w�%����GJ�gkw�h6��v|��l���+9�����yV�  8Mw��OnG�R� `i��0Ro�v��I��v g��`��N��""�����n�k'�f��	 �S(��hG{Q懵S  �3t�;�� ����nDӭ�Ae��/\��?~�v ���`�]���"�K�;xt;��� ��J;�v�r�1��  �Ci#�oD>:��� [J�/�{��-E�s���� �>w�%�I��D�����u����9g�p�; ,��#O�D�G�Y�  ��2=�vt#J�� ��J�^��v�*kR����jw p����3׾s!"���<��M�OqvJ���]p�eQf�ю���ƵS  ���,��F���  W�ߊ��Y�ZK���̗kg p���T?�߈��;xt����sv�fmO2��W�<��ȓ�%��  F�|t'��-�+  <��ƅ�ԩ�AE)�7j7 p�����_��A����<��"��������G�B+%��A��~D;�]  ,�2�D;ڏ2�} �#KM4C��Z�>t�S���3 8=� K����W#��<��a?�&��`����	 �C��Q���(Ӄ���  �]�6��ȓ;�{ �G���H���T�6�?�� ��1pX6ׯ79�?��������N`�M�`��6���ȇ7#���  ��)�q��Q��7 <�f��x���ʿr�S��� �w�%���\�|��@�υ�A�V�x2��  �S"D;ڋh�j�   �,�"���LǵK  �@�f�B�ĭ��R/���� �t�j�lJ���	<��A/�]_r9;9���]��EP�����AD��9  �J(���D>�Qr� ������%w�Sʿ󾗯kg ���� �ȕk���ӵ;x<�]o�lMf�(�s PW9�ڞ��ٓU  ��W�hG�QZ�s  ���ۈ�ݨ�A)]����v� ���;���g�x|����	���Ѽv ��2?�v�wr�  ��6��F�#�  ��f��tkgPA�� xz� K�W������<�a��^�v+��� �(9��v�Û��]  ��ez��fDɵc  SJ�l\��T�����+����kG �t��D��'�;��sqkP;�5p85p��Vf��W�g��S  �u�E;ڏ2��. XH��F3ة�AmJ��v O��`	���>�J\��������N`ŕq4u1 �K��h�7"On��  �W�ȇ7"�. XH���;���9kJ�������� <9w�%�F�������ub�߭������K�� k�D��"��#Z� ��R�юo� . ��h���S;���D���3 xrƒ ��o�?J�z��ŭA����Ѽv ���΢݈r�zD�`  ���i���(s� x��D�q1"R��U�ڋ���Y��'c���R��ED8��.�s�� pfJ�|ty��g�k   �]ɑoD��	� �/uz�۵38G)ť�Y��� <w������(��<�^��́�%p�&� p&��������v
  �c+�q��%�N XM+��P�:i"�Q��'c������K��휃R"�w 8U%G>���fDik�   <�v�h?J�T  wu6.D�N��KJ?|�S��� <>w��������߬�����=���8��#���Rf����I�  ��Q������{�=�����|�{fzf�\�93����J\,[ #C�1ج�����肍��H8B�J>��#�Vk�S�8IU*��W�*c�C�r�J*N�S`�d�����t�t��������sfz�ӗ��/xVmU������ݏ<�. ������t	W%��J� ��;��jZ�xDtJw���;�X]vx��w:py	 &��W���)]  0a9���h�GϾ `���R����\�TUo�y�co,���1p�B�=����Kwp>ۮ�sEzg� pQy�j;  ��u�n�f\: ��ji-R�o��!WMt ��`
���C�T����Z_.���p� .��W����  �Gs��!_ ���V6"R�tW ����o���� �?w�)s��O�*"}O��gu�� s�F�&Fcc< 8W� �������ȥc  �IUTݭ�H�K�d)b)uW�f��;��i7�c���r���rz�z; <0W�  ~G����� Xh�Չj�Z��@��}������ �w�)r��<�PD����OJ[k�\�Ӂ�; <W�  ^@=���n�ڿ7 �+-�FjwKgp�ҵN���� �w�)�j��5ͨ����}�r5��>5uԽW�  ^L����G�K�  S�lDT��\�T���ȣwVJw ��� �����s��/���m�����h���t L�<�G}z7�>+�  0�r4��h��K�  \����n�9ݼ˷����-]���0%R�>��Ϭ*��\3p�j��Ƒ�� /��W�G�j;  ��ʣ^Խo� R��Q�\+��e��co�U:��f�0~�S7#���3lcm)ZU*���蝍J' ��r�  ���aԧw#�� X<�Ӎ�q�p�U)}���|G� ^��;����"b�t�w�?p�:'}?,��h�{���  LB���DJ�  \�jy#��������� �4w��n����H�-���-uZ����-W�ir�������a�  �9�D�?���t ��J)��f��ͳ�7�r�[KW ��|V������������	,���8��Kg �t�ύ-\m  �4yxM�0¿K $U��F�̫���n ���t��O>�W���پf��չ�w� ""�x�����A�  ���ǃ�{�M]: �ʤ�r����\�TUo�y�co,��3p(�i�߈�������R,�}�ruN���	 PV������Gd�
  �+ӌ��ݍ<v� X��zDk�t�"WMn�p�
 ^�E@!�����G�w���b���������; �+�ύ)F��)   �)7�����. �2��fDj����T�m۝W�� �K��T��>�gZ�U�ƪ'��:'�a�\� J�ќ݋�w7���  Xp9�ٽhǥC  �F���nED*]����i�_��/eX	P��w=�D��^����^_���W�����v On�Q��Gv  `��Q/��A�� ,���D��Q:�K�"ߵ7=~�t �g�P@�T?�yׯuK'�`N�� ,�fx��݈�w   �T�Ϣ��G4u� �K�:�H;����u���� ������;?�G#�7���b�V:���*����ǥ3 �j4uԽ��g�"�%@  ��֌����p2 0������S:�	K��K;��o�t ������H-���]��R:�s2�� �!��Q�ލ���S   �_���wy|V� ���hu�"���\Iig����� �.ߴ W�ֻ>��#�7���bڭ*�֖Kg�`���� �s�����("��5   <�&��A4g'�C  .WՊje�t�R�y�k� S���ܹS�\�x�.������T:�s�3p`~�� ��g"��S   ��<<�fp�t
 ��I�H��Jg0A)�C�K�{Kw �,w�+����zOD���\LJ���*��F1�]�`���8��aD�]  0/�u�0"� �ZZ�Զ�+U|�w��`�p~�N��z��X]��N�t���v �Pn�Q��#�z�S   ��YԽ���.] pi��͈�S:�	I)>�6�_� w�+�{X����;�������0_��i4�w#�Q�   .S3z����� ��J)��fD2ÛU�?��[*���|�\�G���D�����;����7Wk8nb0�� ���M4���g�"�k�  B���D;� ̧T��Z�*����*�z������ ������z���_Y������-��:N ����aԧw#��S   �rM4���# �)��"-_+����*�h<z�]�`��\���'�#ҏ����ZU�����,�{=W� �u9��q4���\��  ����0����!  ��ZZ�Զ+�)������� Xd� �������\����hU�t�ir��G�3 ��r3��t?�W:  �)��'��Kg  \�je3���`r��bo�U�`Q�\�{O�"��WJw07�uK'�������\: �%��ќ�G4�  ���M�0"��' 0gR�Vw+"��ͺ*�/�q�u�]�`Q�&�$���fD�����u�be�C�\��ްt <��D�?�fpM�   �T��D8� ̛���VDxK����C���a�p	v������77]o��{� ̘<F}z7�xP:  �YP���GdH �%��"-���ࢪ����{O��Ed�pr���3v.�,�ccu�t�w6�Q�G fE���$��~D�K�   0K�ѳK7��%  U-�E�8�7��P� �+�`�n�}�OD�7��`2v�VK'���N]o`6�f��~��I�   fU����G�G�K  &�Zو�:�3��*�ޝ���Jg ,w�I��ǭ*�GKg0�v[k˥3XP��g� �e�� �����   ��M4���c�? �y���݊Hfz���Zq��j�������_���.��d�l�FJ�+XD��QGu� x	9��q4�ÈhJ�   07�h��ǃ�!  �S���nG���J������� ���`Bv��X���Z�&�U��qm�t����v �Wn�Q��G�J%B�8    IDAT�   0�r4��ȣ~� ��I�NT+�3�����n X$� �R|0"*��d���FUyz�2�z^��tʣ~4��ͨt
   s�� s%u����Jgp^)����~�w�+b�07����#��Kw0UJq�Z�t�w6��.� ϗs4��hGє�  `A4��h�NJg  LL�|-R���gV��q���
����V������ؾ����H�8<9+�  ϓ�qԽ��cW�   �zyxb� ̕je3����|��ƛ��*��� .h�=�xC���;���"v6]o���Sw �G��9ݏhF�S   X`yx��t �d���VD2ݛE�����V��y�[����\����r,w�礌��(F�t D�M�(��QD�n  ��<�E�?��\: ��VTݭ�H�Kx@�J_�}�U�_�`��\�λ>��H��L�Ζ��sx�z; ��zu�n�q�t
   <O������ZKQ�l���R���#��Y)�0���k��RN?]:���X]���N��ᩁ; e�a/��~D3.�   /(�Q�#��; 0�R���Z:��Rz��J��� �����n��}_D���Lέm4R��`�qS:�E�s4��hΎ�<   �^}u��� ��ʵ��r�P���;��o�t��2p8���'�s�/����Ni��PJ�GQ�>y<(�   ��� s"E��Q�K�� R�����/�0���#����Jg09��SR��'� \�<�G�ۏ�u�   xpF� ��HUTݭ�d�7SR�?���ǶKg �#߈ ����^�">P���q��Ҏzg1��� ,���8��QD   0��aԽ����X�ٖ���#�H�S�O)���Z�� �����T��X)����Ni�� X �G}�y�+�   �ь��� 3/���Z�(����⽻o�Э� ������{�[#�w��`r\o��q�Ľ��t "�Ϣ��G4��)   0YF� ��H�n����ܷt�^j�t��1p�_��i�?_:��r���N�"�� ̿��I4}?�  0ǌ��9Q-�GjwKgp�r|����<R:`��ܧ��[��_S���q��i�oP:�y���{��'�K   ��� s��nD��Jgp?R��r��� ����>�r����?V���r���zg�ǥ3 �c�F}z7��N  ��c� ̅��VDj��>��}�m�=�; 慁;�}������;��ۙ'��py�M� "ץS   ��� � UQ�n����K)u����; �o>�������F��P��ɺ��V:��s���Y� �Q����9;��\�   �1r �@��Qu�""�N�e���Ν�?��� ����eT)�|Dx���Z[���v��q�,ƵU ��\��>}&��[B    "�����: 0�R{)�������8w\q� w��pk�w�o)���q����w�z; �G�hz�.�   ӥF�?0r fZ�t#uVKg�2������}��Kw �:w��ʽ���U���L֍�n,w䧬q��q���I����E���   ����^r#w `vU+��+�3xi��T�t��3pxô�x����LN�J���if�ۿ7p(���MԽ�ȣ^�   �~�Y�=#w `�U�͈�R�^R���o��;KW �2w�p��O�*"�p�&kgs5:m_}���q�t s ף�O�F���)   0;�h�Ga� ̮��VD�.�K�Z?���$�9Y���v�~."���#�V;���ǽa��M� f\����G�t
   ̜<<7r �Q��������U����|��Jw �*�p _��;��c��L֭�kQU�t�]������8��Ks   py<x��k �ٔ�vT�툰��Z)}x��.�0�����?n59�|�&k�ӊ��+�3 ��&����3 �U���wy�+]   s!����Kg  �[ju��n���E�7[���Kw �"w�/����O"�Jw0Y]_��e����~d�v8�\��>�Q{P
   &)�z�OKg  �[j�DZ�V:�������ï*�0k��s�;�ܭ"�F�&ku��k˥3 r�ؿ7(��ʣ~4���\�N  �����Ezc 0����H��������~�t��1pxN���ۥ;���o��N���8<=�qݔ� `��hG��"�+@   �25gǑǎ�  ��Zو�^)��I�=7���?P:`��D�����]����Z[���N��������	 ̒�D}�y��   �J�?�<��  8����Z*���j5���� �����;�鉈H�S��*��}��v�C8����t 3"�èO�F4�;   �j�h���k� �*E��Q�K��ER��t���S�; f��;��vww�)�P�������r�U:""����p�M� "ץS   `A5��"7��!  瓪hu�#�i�ɹ�h��� ��b�B���'^�>R���괫��\-�Q79O�x99��Q4���ȥc   `������ 3�jE����)���~���-�0|����ߍ���L��7֣�R�����{��CE ^Bn��D�K�    �����)] p.�Չ���S%ŝ���\mx����}�o�H�Q���Z�vbkm�tDDD��;�� `��z��݈zX:   �b�8��ax� 0�R{)����|���+;�?R�`���{�)�t��ҳ��aZ���h� /,�Ͼ�<{�9   L�zM��t ���N7���|�����<�#�Kw L3w`!���㵥;����.�Kg��p���O��F��   `��� ��q� �s���"-����wm�++?^:`����>�U郥;��v��[[��3�w��G�?�� `��M�0�ٽ�%   �ȣ^4���  �V-_������R������[:`Z��j������L���k�n�Zcz�����MԽ���A�   ���=� 3��nD�Lf�A�Xʭ�S�`ZY����o/��du��q}}�t������ްt S$ף�O�F4��)   �4��ȵ���Y���݊h-�!"R��v���?,�0�܁�q���ZN�o��`�^qc=R*]��i���y4������)   ���h���q� ��Iύܫv�"���g��{�8 �"���H+g="^Q���ھ�k+���;F�&O���g5g'�#"�N   &%7��"rS� �|R��vDj�.YxUJ_��ʯ��� ���X��>�5)�Kw0Y�V__+����q?�# 9G�;�<<)]   \�\G��P; 0êVTݭ0!,/��C;����� �ķ� r���dD8�=g��햯2�G��ؿ�z;����8��݈��t
   p��a4���  �Z��V�""�NYh)��fy�'Kw L����n�ňxo�&k�ۉW�X/����� �N�Y����"r]:   �
�8""R{�p �����Վ<�[wQ)�a�˾���ͯ}�t
�4p��k;{O�N9�T�&�J)^y�Z�x��#>w�+�@Ayԏ�w���)   ��Ó�#o� fWj�D��Y:cѵrg��KG Lw`��T},Gl��`�v�Vc��%$L���A��� ��9;�fp�t
   P@38�\�Jg  �[�D��Q:c����[?�]�; ���;0�v���?���t���Ԏݭ���<9G<}�z;�b���"OJ�    E�h��M]: ����j�����I��>�u?`,<w`.���_��|�t��ʛ�R�
x���AG~� X8���wy�/]   L�\G�?|�*
 �����#-���XX)�Wvn=^��4w`.����L�*��d�����J�t<��� �)7�{���t
   0M�Q4���  R-_����XX)������#�; J2p���'�`�齥;��N����{B��sp2�3��J���G4��)   ���A4g'�3  .�Zٌ�^)���R�V���� %����;�&�"�U:��z���hU�t<��� �'����"rS:   �byxy�/� p!Uw3��\:c!�������� ��s���ΏF�ז�`�6V�bs�LL���3��Hsv��+�s�   `4�����t ��hu�"�N�E�r��swl<�����;���W�>\���jU)^q�Z��9G|��t W"G�?�<�jq   �A�h��� ̶����m�^BJo�~��Jg �`�̉�R����n�&����u��q�`A�&��A�W�   ��{�p �LKճ#��*]�p������m�� �j��\�y�'�7R~S�&�Zw)n\[)�/���^� .Yn�Q�ލ���S   �Y֌���  ��TEk�����K����/]p�|� 3���<u3�濍���-LN�J񚇶�U��)�%O���K� �,����"�+�  �	h�)Ej-�. 8�TEj/G�j�R�˯���~���ߗ.�*.�3oT�����;��WܼKm_SL����0��xM߸   ��|v/���t ��������d�qURJ����xD�	,�2�L��{�m)�ݥ;��͵��^_.�/���,�q� .I�����#   �eh�G��� ̶T���n�_���7�x�G��� W�70��SO��*=Q���j��xō����r�����3 �$��8����   �\k�}�>{� �m��yv�n�x�~�ڛ�Q:�*�vfָ��D�xm�&�7ף����tz��Q]:�����#�z�C   �EЌ����  ����D���t�bHi��j��� W�U: �<n����9����\�Z_���k�3��M���q4�� ̗�<��r}V�   X$��c*��T8 �bRՊ��D���*�*�q��������v���d
̜�x�/,�����\鴪xō���>wԋqݔ� `��:��~D=,]   ,�<<�<��  ���^���.�_�VT��wl?���C�9����Z�x}�&�;ע���t����a�t ��QԽ�͸t
   ����qd�> ́�^yn�ΥK���o��� ��#S�L��{�kSJ�kDtJ�09ׯ�īv��΀��gN�;����a4�È�f   `
T�h�ވH~� f_���Θ{9�3æ������.�p��fǣw�)�/�q�\鴫x��z�xQ�a�����E����q;   05�� 07R���F錹�R�\��?]���3cww�F�7��`rR�x��F�*I�^�=8��KW 0	���s?�`   �K����  ����i�Z����?�͏K���`�̄��|����L���j�w�gz��FqxzV:����#OJ�    ��|v/�ؿI �ZZ3r�t�ʭ��bo�U�`�܁���v�_����)L��J'nm��΀���}�r f^�Q�#�z�K    ^V38�h��  a�~R���G_��Kg L��;0�n��~0����;��V��ջ�R�xqǽa��G�3 ���D�?��]>   fDn��F�\� `"�ܯ@��k7����Kg L��;0�n���刏��`�^�s-�ھ��^9��0�ru� ��.   x0�(��q�
 ��1r�\)�ͦ���Kw L�u!0��ܩZ��#b�t
�sc��k˥3�%=s܏�p\:�s��8�ӻ�7q    �)���b 懑��J)��ƛ?��� �b�L���������L��R;��V:^Ҹn���^� �)ףhz��.�   p!��$r�~ `~�_��������! ��* �Bn���_���/#�S��ɨR��<�Km_=L�O���� �(��hz�єN   ��<F��F�T: `"Rk�������S�O���kۣ����_-�pQ.���Ν�ʭ���)L��7ף��.�/�?���~� �!���¸   �+����t	 �ĸ�~yRj��[~�u�; .���:;���_���t����7���΀���'��F 0s��z  �yU�9;-] 0Q��Z�����'�J��'Kg \T�t ����'����X*��dt�U���fT�Wg2�N��sG��̚��$��^�   ��U#�:�*o� �Gj?7��eC�MJ�t_��?���_�?J� ����ɩn�/G��3�DJ��ڈv��ӭir|f��t �9�y��   X��(��Kg  LT��i�Z��Su>����� 8/�C`j����_N�t�����X]�΀���Q/F�t �-G�?�<�jn   `��&��aDΥK  &�ZZ3r�����r��\���j� �����O�6W鿊���-L���r<|�1~��٨��z�^�9 `F������t	   ���MDΑ�˥K  &*��"R����S�GJ_���?�/{�����t
��r�(�Ν*W�#�zN,wZ��O�2>��k7 �!7Q�"��%    ��Q/�_: `⪥��V6Kg̓�T�/�z��J� <(w������#�)��dT)�#�6�U��)�N��8:5��	���w�j   @D4�����t �ĥN��}�R�׌�ʏ�� xPև@Q��>�����ˈX)��d|٭��Z�ZL�_����b0�N��|~����   �wT�h�ވH~� �O�E�7�_T�yT�?��?����t��r�(��;��?
���qs�k�����Qϸ`4uԧw��   �X3�fp\� �R���s��=�wQ)�N^j�b��J� �/w���[��)}}�&cu�__/���lT�gz�3 x�G�ۏ�u�   �����ȣ~� �K�:+Qu��'"�7^?�=?T:�~����y��oLM�_"�S���k����WlG��)f�o|�(����3 x	�E�?��M�   �)WE�v=R�. p)��,��aD��)�-�ɸi�p�O�ߔNx9���������rj���s!��W�^3ngf���L9�v   ��D�?��_ �|J�娺����Xo���� ���r���?_]��ɸ��׺K�3ྌ�&>�Z:�����hz��    �Esv�t ��I�%#�	HU�7������ x9>�+����o�����h�n��6V��5�7Kg�}�wO���Y� ^��K   \L����R: ���zM�0"K:�����W��GJ� �܁+��zj5���q�\X��ջ�3����� S,���    ��#7��  �&���Z�
���K)=�Zk�L����S�2�n�3��+Kwpq�*�#�6�Uy��nr|��f�Vyԏf`�   pqM4����, �<{v��痪���x�c�Z������ĭ�'�5"�W���x��Ft�ڥ3�}��I��^O0���i4���    �E3p� �o��1r��V�:�x�-X+�B|����������?�������X]*���^���3 x��4�[   &-�z�G�m �o�3rOf��Rz͸Z��� /�';p�:���GīKwpq�k�qk{�tܷ���[�3��F��    ��9;�h��  �*�:Qu���-U��~���t��\�[������[���[Yjǫw��΀��'17�3 �"��    W 7Q�#"�. �TF��J���{�7��n��/��4����ݜ�S�;��v��GnmDU��)p�������W�Msvb�   pU�Q4g'�+  .�����*^��X��; ��Os�������V�.&��/�݈�N�t
ܷ���[�3��6��I�T   �R�F���  �t�Չj�zD�qyP��~h�͏S���3p.��>���'Jwpq]_��n�t<�O}�^��M� ��q;   @9��(��Kg  \�T��Z�6rp��j��x��\: "§80q��z��#��&"�J�p1��V���k�3�����Ӈ�� |�fpytZ:   `����8��JD��1  �*�*R{9�x�t��Hig�Y������t
���d=z�M�_D�z�.fu���y�t���z    IDAT<��Q���:0�4yv���#   ���a4g�  ���K��#���HU���?��ו� ��L���ΏE�o(���tZU<rk#�̐�#~��{Q7�����    �%O"���3  �D��Qu��L�����fi���;��-�b��L��w��#�c�;��*�x��Ftھ"�-O��w6*��s��   �S38��M� �+�Z��V��D��k�/�>T�Xl���|���?��Ɲ��[��W�n���R�x ��Q����� �9��(�_:   ��#�:Rg�t ��HU+R�y4(�23RT߸������??]�XLK&"���\D|U�.���jl�/�΀�49~��{�s� ">�ݸ   `������  %����nGD*�2R�T��{{�(E������"�_(���l�-������>u�$�Fu� ����^�    �C38�܌Kg  \��^���F����?�}��)�,&���������&�����]����.��+ڊ���l9:=����� �q;   �L�:�Z�� �"��A4���������������O���)�bq���&�1��gZ�U�#�6�ۙ9�q�z�t a�   0��Q4g�� X,����F�ِ����"�ؚWʇpn�����Gķ�����������u����3�b\7�3 ^svb�   0���4�xX: �J�N7�e#���R���>P�X,���r��xmn���J�p~��ڈ͵����>wԏO�uQ����$���1   ��K�h�݈H�" ���F>�W:c��<h��?x�?���]:X�:ܣwڹ�%��g�C�׌ۙI��Q|fߘ�4�v   �9��hǥ+  �\��ii�t��Ki�j-��x�N�t
�܁����c�Kwp~[k˱��Z:ظn��~�8r.]�،�   �O"���3  �\���cG��u�;�GJg �!� f��;������#�U���Y[�ė?��7 3�7>s���� ͸   `�UQ�]�T9�	 ,��y<(�1�r�0��|����V��o.��m{�͈�+a�>�:�*��a��L��Aϸ��fxj�   0ךh�G�U� �⩺����S-E,E��y��J�`����S՟��GJwp>�*�knoF�壟�s��gOKg ,�fx��^�    .[3��̿� �(E���Z*2�R�}���(��7+G���=�ݑ�Jwp>)E�zw#�K^'�����ͧ�#;PL���   H�D{�* ���s#���楤����o~�[Jw ���xY��>��H��;8�����ƪ�K�=9G���cT7�S V��9;.�   �kGٿ� (U��nG�V�i�j��_�y�}�C��d���G�s�~%"6J�p>77����-����N�?*����x���   `!�ڿ ��jE���L,_L���z���*��'���Kڽ���H�Kwp>�K��uJ2��{�x��W:`a��0��QD��)    �ǃȣ~� �"RՎ��f�/.�Z߿����x�`������}����yDx���.��+ڊ��Q������~� ƵW����Q4����9   @���HU�t @y|M�0�za9ǧ���~��[����"�m�=��%��gR�U�knm�3�r��w�=6n(ĸ   ��k�� Xh����f錩�R�������;��b���N?��������yh3:m�̦߾{��Q�����q4}�v    �H3���t @1��i�Z��UU���������~���;?��"ҟ-���K)��nmDw�+"�M'gq��_:`!�f����l�   ����y�egy���s�]��Y�Ui�R��W��Y�L��a��,a���V�m���{:c��nT	am6H�3��тl�D0ƍ��``P-��\n.w?�3��T��*U��y����`��D��y�x<o��3�  �ޕ�d���ye�ŽS?���! 6��fz��;$�݁�ٶePC�R�`]j͎:�; zS�n�b�       �\�Q��c�   D��Ii9vF>��:���� 6�4v ��=W�M�]�Sp���55�)Qt�v'���%e�/�`�yPVg�      g���.+0�  z�))��;-nF~f�C��_�P}�}_��������MMM��L/�݁s7:P���@�`]ܥ�/��� l8�j�R��.     @��v��@  @�2S�?&���PR��#/{��3 t7�H�&߰�j�~?v��@_Q�N�� ��+Zk�cg @�qx��g0      �MhT�X
  z�%J*�b���l�P(��fg9 `�x� ����2�)i,v�M��j�����N��D���K�� Ѓ\Y}I
l�     �z��AV�  �%�,-�;��)�c��������B� ݉�C@�s+��.�]�sSH�Q!�Q���h���j� �I�^��f�      t1o��  =�
%%}ñ3�)I�>����0v���w��M�N��Lo�݁s��i�̈�˅�)���:A�T��N����N=v      6�ZJ�ɸm  �.K��\�ڱSrŤ��=t�~�v蟹Z�9a�/�æg��cn���8w�Li��;X�\��U��B� �9��"o�bg      `���X�]  ]R�*�3r'1ە����@�a�;У���JwI6��fۖAmꋝ�ۃ�W�Z��2 l4o����      �lBG��o.  �]V,˳��Y�\1K~�rŋ�Q������{���Q���n?��fr���N{�{[�ii�; z���
M6i     ���)0�  z�)��J���3�yq����e+��ƀ;Ѓ�g�^'�Wbw�܌��m�`�`ݪkM]\�� =�;M��     ��5��#   �DI���<�i*���o�3 t�
=frv�.�}FR9v��@_Qۧ�ef�S�u��::tlY�K ��x�V�/I�     ��3�L��b�   De��҂�ӈ��+f��|�����|9v����K���h��K����W*��>=�$a�ݩ�:��,0\	 �CG��()�N     @���<tbg   Dg���<;#w�$y������� �pz��R��^�g��&�|fD���5�S��G��jg�S ���L��(9��      �H�P��  ��4 +Tbg䋩b���u�o�c� �7&&�1yݾkM���8{��v��\Lc� ����՚�� �[<(�-��      �h���\�]  �IeXJ��3r�L��F�0v�|cj�[fo�(��4�g�L�ljXC�R�`ݾ7��ŕF� �-��j��s4      "�ڲBY�0�   z�))�坦���Q��v^uom���b� �'6����-i"�����)8{۶jd��xн�W:Y��� ����R��      ��
���  ���J*��,vI���ҏ��~�h� �Ā;��M���ʹ;v���X�&�+�3�u[�����+�3 ������bg       ���Bs5v  @.XZT�7;#W�첤o�C�; �������]m�G�a��1:X��C�3�u�5;:x�*g! l��\��k�3      ��emY�$KM   ��(ɥ��af?ҷ�꣍���J� �§H`�y㾱B���c���V��>="�6"t�V'���%e��v �Hު�[l�     @>y����/^�  HV(K�s�$I&���/��q���c� ��:�T����uY����R��vt�,������) �S��Ph.��       ��g
͕�   ���KI!vF~���P����s}�S ���&4yݾߐ���8;�b��gF�&L��;�K_V���b �H�����      ���vM��bg   �%J*�b|�Qfz�J��G�; �G; ��5}�M?*�-���[��
i��gFU.�8F������V��3 ��x�(�%y�      �x����/�4  ��Y��;��)���?ٿ�%_���۱S �� `���?�H��n��K̴cfX}%��ѽ�/�4�\�� �ŃBmQ��      8{�)�VcW   ��d���9�[�����]�@|����?`�����3�.�R�E��^��MYX�� ��]YmQ�,v	      pμ�&�Z�3   r#)Ji)vFn�i�B�1i��V��� 6��=7���bw��\41���r�`ݖk-}��r� �1���$�v�      `�B�*���   �	SZ�,��������� ��lS�ݼ��N�]`fl@�#����՚m<��w� ��B�*e��      �3t��x�	   I2��%y��$?,��rً����) �`�;�����}B�p�<��>M���� ֭��t���� ��BsE��-      l�Z�g��   �aiQIy(vFn�TR�����<�@�]n���K������/��	~E�jw��YR'�S ��x�.o���       ΫP���b  e�~Y�;#7�l{Z��@i�  �79���&��$�݂��_.j�̈���U�NYp�?RU���N��❖B�;      � N�[��   ?,-�;-�Y>(I2�������_b� �XLZ]j��dZY�k�fb�੕��vmU!��t�\�V��h�N���Y[��(�/�      �y%�㲴;   7<t��{��[6o<�����v� �iK���%����WL]���vt/w��+��F�P__Z     `���   �$YRPR���'�A�O�������0q	t���z������SKӎ�#*xԢ{=trEյf� �-��j��g�K      ��3��j�
  �\�BYV���f���l�=�; l�4v �s3��?%�G��\3�v̌j��;X���_n�� ����KRh�      6N֖J��  �GX�$��,�z�%���w��_������- .<d�.23��IS��
�[��.��`��vt�պNT�3 ��Ɗ�qs      zO�W%��   9bJ�F$c��O\韌���c� ��x�]�-�%]�OmۖA��cg 붰���y���Zk�v-v      �g
-�O   �&I��Ǯ�3mI��I]y=�G�M����.19;�V3�z�<���~M���� ֭���wO��� ���톼�;      �+k�
%Y�(  �#,)H�Ў��vq��������b� �p�Tt��7|��}L�����`YO�� �m��ҡc���	 ̳�B})v      �����*�,v
  @nX�$�N�C�$/�u��j�����- .�$v ��6��}c�ɧ$q�J�V��t��н�m:�p; l4����y       ���Qh�Ů   �SR#���$(���+�~I� O; ���m��\��.�����1="c��T�����U��`cy85�Ζ      �4�Z�g��   �bIAI���0ӄ��S�=W����Kc xrS{��W�~#v�\��j�̨
)�Нꭎ]Vn�����KR�%      �D<�()U$�e
  ��N-��=�$�L��%�bc��w�np~1�����M�w����in�D�ό�\�o�S������:��`��Ɗ�i��       �˃d�,-�.  �+��7E?̒�ŕ�/�r}�}��np��rȡ�׽w4�R���Tb�3��+1܎����?��6�� ��BkMޮ��       rϛ��Љ�  �3��2"�?�/���щ��e[� �O8 w�J��G$�]�'f&m�V�;X��#����`�y�)o���       ��+4�cG   �%%}C�3�dƓ�'�9fb�M���@�L_7�f���O��!��cg ���N���Y� �9���K�<v
      �=<�Y"KY>  �X���9����ʎ������) �9܁�x����R�l����M�Tbg �ׁ�U5Z����P[���      ��򬭤�'9  �
%y�!�l�bI���W}�����[ <3|�rb�u�M<|JR)v�ؖኦF�cg ����Ѫ�MN���se�%�9`      �OP֨Ǝ   �K��ĮȓTI��&w��L� ��@N�J�?����xb�e]<1;X������F;v
 ��P�JY+v      �ݲ��]�]  �;V(Ɋ,�|���f��Ǥ9�c�.�0�����I��݁'6X)�ҩ������:x��v �%4W�F�      `S��C�  ��I����;#7,I^6~Mg.v��Kc �n��=ۂn�T�݂��+t��Q%��N��#��u�� �4����      �&�R�dž�!   9c�B�o��^�w��������np���D49�wP�n��709T*��|fD)���B�@\�����      ����&  <K
��`�<I-)�����.���1�Dd��,�Y�;�x�4ю�<&�}Bp:��p; ��A��$�c�       �Rh,Kbg   �NR��r��0ӄ�'u����- ���@$S�7��\o�݁�K̴cfX}�4v
p�ܥ�/k�ފ� =ʕ�%�b�       ����J�
  �\J+#�1�3�h|b�{bw 87LoLϾ��dv�$N�匙�cfD�}��)�9s��j��p; ���R֌�      l~�#K����   _�dI*�4b��Y����/�F��}ߌ���pL�`��{�$�H��n��]<1��
���>�@|��*��cg       =#4�O�$  �i��'+2��(OT(~x�oyV� g�w`���M����;�x۶j|�/vp�n���Ӑ�Vcg       ��3��J�
  �\J�Ò��3r��F�ʟھ{�1�0�l��={���_�݁Ǜ�hr�S��>�@|:
���      @O�vM��  �q̔�Į�3{�r���� ��s�2}�M?��_I*�n��F˺dr(vp�ܥ�/3� 1yP�-H
�K      ���Y[I�"�b�   �%��A
��)�a��D������k�[ <96�`���h ��"�?vN7T)������9{ds{u�; z�+�/I��      z[�(4�bW   �RR��]ȧI����mύ���1�l o�3�bw�t�墶O�X�.��v ȇ�X���      �o��36�  <����H�|1H���W�e(v
�'ƀ;p�M^��W%�J���TL�}zXI�t;�K��G�� �y�&o�bg       �>Wh,ǎ   �%KK�b�\1�g���ͱ; <1� .����Gd�I*�n���i�]��T*p��%��cU���> 1y��Ш��       p&2Kd)�g  �diI�nH��)�af?ַ�%��~9v��1�\ ���ѾV�}V�%�[�41��:���?t�,��j��p; �䡣P__�       ��Y[I�O2�]  ��L���z�\��~�o�U��8p�wc� x���^�����x��t����˅�)�9yd���d� �rW�W%�K       <����;   �,-Ɋ��3�Ŭli�S��w&v
�G1�\ �����~5vNw�԰�*���9iw��?��p; �@hT���      Ƚ�)o7bW   �RR��>��]��ʟ��l��)�0����?x��?#���ڶeP[��bg ��	:p��F�; z^h��۵�       Βg-%�ʩk�  �(3YZ���Kr���_/���{w� ����7}�����tY�<jz�_ӣ\������?��f;�� =�;-y�;      �9qɃ��,  �3Y�J���LI���]W������f���%��ͤVk�O�scw�QcC}�����G��[�@t:
���       ���uy�;   ���d�H>�'.�ȖW���.z��y2��=����x�pI�L�� �I�����-2� y�P���\       �+�FUr�܂��    IDAT�  �?fJ�FbW䎙�x���mW^���e������]&���x�@_Q�M�,v	p�ꭎYR;c� � 4�\�      t;�Zk�+   r�
%Y�;#w��9�-S7�� z�K �Юk�Wn��K������.�:�4��G�������0� ����v-v      ��!k�
eY  ���P��뒸��4�=�|�����|9v
Ћ�������{%���8��&�|�
������:p��p; �w���j�       �+4���  ��DIy(vE.��������@/bx&g��{�~-vNIӎ�#*x��{,�Z:x��,��* 䁇�B�;      ���
-nm  x"V�Hi9vF���--|jr����NzS��:M]w�N3���8%1ӎ�UJ��)�Y[\m�б��3� ����p;7j       ��7פ���   ȥ�oX��>��]��ʟ��l��%���q��ŁFv��]�S �I�Mk��;8k'�u=tr%v �1B�*e��       .��LI�;   ,�L�3}�؎��x���޻c� ���6�:L/e�U�cw������t��K5�_�� x��\�w�3       \hYSޮǮ   ȥ�4 %�����2~��_;���hj���s�?���)�c��a�����UYX�� x�4�-      �"4W$�3   r)�֩U�8�'��O&~� v	�p���ٛ/��������`Y3c�3���.}�ĊNT� �2�F5v      ����Ԑ;   �Ң��;#��l����Uo��lv�g�����|R�x�H���.����w����ZXi�N �ƕ՗��      � o��V�  �\JJ����3�)��
.����Y�Z
��E�; U����+�@��G�ZZk�N �!4��Ў�       �Ш��T  �ә)�cI��I��붼�mo��lf�����W��}��Ut�b��3�*���A�u���ǖ��`x �&��䭵�       �rI&+�b�   �%)tN���%�Kv^����{�;،�����^���L�GWH�Q�������?R��� �;������       r�[k��9   O�ʃbl�I�!)||�+~�c� �S��S�=W(�KI[b����L;f��W��	�_���;��hq� rǃB}I�63      �+4�cG   �%Yi vFn�4����&w��`�`�a�x
S�S�tU�^g&]:5��r1v
�jͶ�YR�b�  Ǖ՗$�b�       ȓЖ�j�+   r))HI!vF~��p�7�gb�=p^�<��=|�)|F��Dw�Ġ&�+�3���Ro�c��[� �BcY��%  F��
mI5I2�%%g��������5%�oX& �X������_�36��~�J��~;���6� ��)Q:8!{  �䝖B}!vF���y���|w�`�`px�?�����W%M�n�u3c�돝<��զ�{bY�l; 䒷�
�j�  �œ�[X6%K.���$�%�]Z���J�!IZ�aɃ�]V��jAi�^Ȫ#}�k���� ���?�T��N:�QV�'#&��+n�h�y93�4fҘLcrui�d#.3ٰ�c�o �+�)����   ȥP_�w�3�����y��+v
�0��i�\ajr�d�:vJ���%�,�A����ux~5v �Ix�V�-H� `ssi�d�.7�1�N(�{fvL�*�L��|���+�͝�� ��q���ƉN1Y{�y6i�)w�V���t��ɦ]���㱋 �-���
}�3   �ǃ�Փ�B��r�ɠ��nס�-@�c�8��}7�����n�����#2�Rȹ#k:�T�� x2���K��. `��VevD҃���a)��+U��!I/t��ֹV�T  ���+���&��R�m!hZ
�}���%]*�m�"� ��R��E%  ��֚��;#�<����<~��|��"���ӳ7����))������E��:�$���r�:����^�<�< @wH�2=(��ؑ�:li��=ܯ4yh�o~��� �l&w��`(�\li�d�\�,��]��̴M�+ ��e�~%}ñ3   rȕ�-H�;$��çn�l���1=
<l��oޚ��I�����J�T����XHb� O*�Ǘ�\c9" ��  ���q�C&�����w��3�yr�u���  ���\i�Y����g��]��v��s],�B�D ����o����   �㝖B}!vF�y��;w��Ǳ;�nŀ; Iss�ԿM�!�e�SzY1M�sۨ�E�� �:Y���˪59�
 y�YK��(�c�  zG��a�0�C�:`��{'�N�������� �yr��ŉ��;���.�.�|�d����T�� 8��ҁq1V  �xܤ}\W�gn��S�n�'1@��}�g�;cw���L;������W����Ѫ��,v
 �xP�6/9�k �qj����f�M3�F�?b  ��?�n�~N�G-�+�Y�@w���@�  ��	����b��Ss�ɠ��nס�-@�a�=o溽�n_��du$fҎ�UJ�S�'Ukvt�hU�,�N <%WV[��V� @�{�A��b�����j��  @���+M����9���g��/� �L����p5  ��BsU�Z����_�TW�z�K�eIppGO��y�h�W%����.���P_��I��[z�ز���S Ȼ�\���bg  �N��oX���ۿ��_m�������f�2  ����}���ҳ��?��Bx�����c� �����Ů   ��S[ܹY�����w����t��Ӧ���	�����m��h��I-�4���9�� �{�i*�cg  ��˾���%%�ݼ����?�&�� ��{�ܥ�`/�ܟ��?.�g�tI�. �UIߨ���.  �3y��Ш���
��y�w���;�n��;z��u�����$vG/��%�C�3�'ul����l�nࡣ�� )�N �K�����kf��e�/����Gbw  ����s���n��ܟ���0� ���%�K   r'�-HY+vF��7-�\s��;���'M���WX�E�`�^5�_���O!䐻���-�4b�  Ί+[[�B;v  &�U��%ٗ����N�>�� �f7��Ǌ޼*H?���+M�� ��+J�Fbg   �gm��|���~"k��-���N��R��]׾��<T�$=7vK��/�s눒�G�'�Ǘ�\�d) t�Ш���� ���ɒ2}݃��*��_��Wy  ��7���K�n~����ҳM^�� �AR�x�  ��w�� �W���K}~�͛�S`�=g����w����W�����6�B��}ȟv'�౪��N� �Y�v]�Q�� ��\���If_��|�oh�������  �,l{�\+�<d/���K���cw@WJ
J��Q  �3xP�zR{hΆ{�������;�<�Sz���W'������(��v]4�R��v�O�����%�;�� ��CGam^��N �o�<(ӗ/�kI��?�֯�N  �L�^3wi���d/q�J��� Ί���cg   �Nh�ɛ+�3�F��K�}��cw y�U�[fo�(5���-�[zQb���F�_.�Ng��֡c��d�@�pWV���n �&�ɒ��I��J��<��sGcG  ���kn�j��KB�%��?�L��] �O�d`�,�'  ����w�b�t�f�+����)@1���0{K:m'�v饱Sz��t�԰FʱS��YZk��W�� �MB�*��cg  �íᲯ*���랅��-��  ���^���������̮�gϕ�/��iIi�x�
  ���v]�Q���5��{I�|�ɻ�s8v�7��'L��?K>��W]41���J��qNT�:<�; p��R �N&%�&��f��o`��n�mN)  t�+�/�O^����J�Z�/`�;�^��Ȋ�  8S�6/�v쌮�!|i�o��7nm�n�wlz�o�w����4vK/�������iܥ�ͯj~�� �6:
k�y r�%}K�|�e��V�s��{+'�   6��W�8V���]����S�_!�;�9���	ɒ�!   �❖B}!vFw	�����bg y�M��F_���R��5�.��ҋFʺlz8vp�,��j��IQ �:��j�R��. ����%_0�}��/���?�	   g��z��r��=�ԤKb7�F�B���h�  ��	�%y�;��d
����w�?v��cS�ڳ��%����h����gF�$<f��v��G�j���) �u����� �%_P��QP��c�{b7   ?&^��j\+�W��jIC�� �BI*c�B9v  @�����d���jd!�f�����ش�����r��������6�B�u|ȏZ��CG���B� �:x��Ш�� ��f�w��Lw�Н�u�;	   ]`��t|�[�W~�\���w� 6K�LHƣ  �BcYޮ���.�'2���t���Nb�6����GB����J�^SH��6�r1��|_u����(��N �é���x��FrْI���n/�o�{0v   ����fB�W������4�	 �)+()sY  �i<([=)�e����W�'����W>�� �4ܱ�l�G�jk���ٱ[zMb�˷�h��;��պϯ��  ����ڼ:�K �X���>o�;O;|���v�*   lb�lw��J��J�OH��� �RҿE��  �BsU�bn�\��O/���=bz��t���w�\����E�Mkt�;�$�Kߛ_��r=v
 ����ó .�U�>oJ�6��o��9w<v   z��57l���:��Ƥ�R�^ �#)*c   ��l��Y쒮�����]�;�X�d�Mej�M���ӱ;zѶ-���{f�C\[�J�; �x��Ш�� �M�e�͒��mk~ۡ��5b7   g�x��+�ե���n�Y�gb7�ӱ��@�  �\��e:���;��w�C�pǦ1�����}M�x�^3>ԧK&�bg ��V'�б���N� �3ࡣ�6/n\��Ē��u���f����$�  ��2y��x��u&��W��� r)Q:�EJ��!   9�����,Ϲri�ڍ��=ߌ�l4����{�055�yIW�N�5��%m���4A�5�:tlY�,�N <��j|� ψ��f�l��}'M>Y���N   Η�k�pgG�k��j�_j�b�& �����,v  @�x���X��ѕ<��<;����}�5��)��bS���w���cw���RA���*Mx� �����{|E�YD	 �.ԫ�N=v t�5)�Kf����ٹ��A   ��6���J��s���f����	 ��QY�/v  @����ގ�ѕ<��-ܑ�V�c�'zS��z��^����=o��&�uјJ�$v
��K5YX�� 8�]Whp� �^�,�=f�gTX�������E   @,�^3���� ߣ�_)���M z�%J&$�]*  �#��T�/���^�λ��z�[cg �wt�m�p�D'˾.i[�^��i�����q�K�X��j3v
 �<��QX���m �<�*�]�양0����7��   8�ų\i�V~6��(�R����X�_I�  ���jR֊�ѥ,X��K'�z�_�.6��bn��7���~6vI��tjXc����q�,�бe�5�� 6we�y)tb� @.�4o��7%�>y��g���0   p�~d��������N纠ε&��n��ʸ�P��  ���j�3��k5�~�������)��ƀ;���u{]n{cw�����폝�Wout�hU�N�� 8OB�*��cg @�$'$}&M��:���t�,v   �����81��Zwͺ�W�4;	�&��l�   �
�%y�;�k���V��`���r<vp!�)
]i�u{(s���@cC}�tr(vz�J���-+; p�x��Ш�� ��XQ�ܑ�n9���[縧   �PfoI��|s����N惱� l>VTR��  �����3��{�o�����_lf���\sqr)��Iϋ��K��ڹuT�S���udaU�l; l�������@s5]vo�$�������Vc'   ����?�4k+?�{�z�<Tb7�,L��YR�  ���}���w��k�3��QUt��=7�[����%�b�+����&�SУܥ�ͯj~�_l`SqWV��B'v	 Đ��K�%�Z�O.~�\e   ��ȫo+zkO�ߛ�[�L�xfҒ����   ��"��#s������}�;��wt��7�ڂ�QR��W��i�QUJ|w�8:Y�Ǘ�Z�F �l8���X��/���,K���o?�   �S����MwJ�_0�/J~�x�
`���Y��!   ��v-vFwsoZֹ��]7~!v
p�������;Z*��.���-��L�13��J)v
zT�����U�;!v
 �<�v]���b =��[�}"K
[��� v   ���|퍻B��&){����{ t�D���dܚ   I
����b��3v4��/X�ܻ��O��kL��/$����䢉AM�E q,�Zz�����/� �ٜ�nnA� l^�Z�ܦ`�m���|w�    �����A鯺�M>�@w�B���h�  ��`��y����_r�+�/&6������%I���K&F*�h�`���c�5]\�� � \�ڂڱC �sYK�{�`��蓺u��	   ����������kC���ט��	@�%�1Y�;   ��~޸�O/���=�/&6	ܑ{�?�������pi,vK����cfD�,�C�Z\i�N \ ���9%�*��L���۷�]    ����M;�%����?�@NY�t`B��  8�w��O�:o[��7�� �>1!����oL�m�ݱSzE���m�*�I���v'�бe՚l����;M��b� 8_�I�-^�n^���;   @�L�v�ٝ�~I���E�{ ������   ����O�e�ם������)ܑk�{��ͥbw�41��6�J�;=����б�ڝ; p��LYm^r�� ��[Cf��>|�~���x�   xj���[��|����5f*�N�I�Y�#  @b�����/:y�{��x&pGnM��21}I⋾��cfD�����1��M=tbE�9�	 �YV[��V� X'��u:������w�v�������>gf�,�d&3	��e�E�Z��E�UB�~��o��V��ʖ���u�%��m?�E��@2@��E��~j]Z�X�Q ��9���}]�bo�@�Lf�u���/x�29ɼ��u��+
�5    Z�ș���%���A1k����*�c   b���!�WL�<o�맭[���I	M�Wv��g�#���[:�!C}��@��3Y���y� �2�9�ڜu ,Ԭ��>F��x����   �^֞��E
�Q:G
9� 6\��|W�u  @S`��Ҋ!�(ޖ�#q#1Z�hJ��n����k��)��u�U�� !D�d|V��U� �2�iM�T�� ��?���|��ى�>2k]   ���yɇW']�W�^�ú�Js�}�r>c  `�-�K/M?\��CXg ���;�����/�YRb��	r�sȠ����j=Ճ{fT�5�S  �-��)��% ���w�s�S7�k]   �3����S�Կ9J���{ ���[I��
  ������B��_S���/Y� �D+�ʡgo�m���I:κ�d�cTw��X��3�F��7 �	ByJ�Q�� �'Ⴂ����3}�˺!_�.    I:|�'rչ�פQov.<O|��=߳Z.���   ����5B����?�S���e�ʺMۮ��;�;:�sү�T.k��Q��葉YE~����e�ʴu <?�\����щ��m]    �3�!���8*��)Z� X&�+�[+9o]  `.T��e댶�oM�i�    IDAT��g���ɢup�pG��x�o8�&���p��~�]� ,��ݓ��;��A �)bh(�ĩz ��� J�����Go���)   ��r��O��噍J�;��k�= �����s��3   ����y�:���n/ޚ� �up pGSX�����j�H:ں�������� �4衽3�+׭S  +&*�/J��4�y9�JuU����c    `)�q��oSԫ��6#�����L�u  ��P�RlT�3�O�+
�_z�up pGS�t��R|�uG'����C���c�Uj��3�Z=�N ��P�Q����(w��P��ٛ��    ЖV�uŚ$T�षI�X� K�%J��%ǥ�  ��Ŵ�P*Xg�!b�����ɺx*�������~W.�&�>.�L�u�akԕ���l�����(�: ��b��P��� СbT�9w�sn���-;$�/�    :��[_,ޥ�3�bƺ��l�|�*�   siiRJ���'j���o���߭S��a�����]]=?����-��WY��\�u�\a��G&f'��R����u	�N�^9��WO�v�.�    �4x�����.)��)Y� X�;,�d�3   L��}���'���i���0�S��n�+E�κ�2ԧ��^����G
s*̔�S  �RQJk� :���s��yݐ�     �G�0�3ۯM1�yN�4� �3J���H  �t|�|b�o�l��l�CS�if֝{����o����z������3��i�C{g4W�[�  ��bm�:@�Qu'���?1~k��=    �
��������+��2I�u������3   L�FM�\��h_�]^�m�E��a�&�lܾ:��J:̺��e3^��F��[��MU��=�j=�N �iM�� �+J'��i�'�n�?h�    �h���#\��+Ʒ8�A� O����%Y�   S�|A
,�\.�PM�˿d]�2�abݦm��қ�;ڝwNG:���u
��l�����(�: `!�}/"�� ,������$�ţ7�K�9    �=;�[N�z�yR<κ�~$]Jz��+   L�FE�<e�Ѿ��o�������:�E�cŭ�x��D�����F44�c��6U��葉YEf��c��b�b���������;�X�    @;>c��»��ARb���|�*��^�   S�����쾆�={zǇ'�C��ƀ1V���k��s?�t�uK����F�3Іb���Uq��F �d�VR��Xg h'��ɹ����۳���s    �����'(T�/�s���$��x%}Ò�
  �\|?��b�;��]z��Xw���V���g}\r/��hw�]%�8Â�B�C{g45_�N ���p ���K���tm����/���U6C    �
+�s�D��;o8�	!�]�'ȩϺ�$EŐ�gs�!   f��(�˒��^.ι�z���^��k�l�Hlp�
�x����7$y�v�x��RW�?f,�z#�=�*W�� :[T:_�B�:@���sɧ'���uC�f    ���^���uo���V�Z� �|Ϡ\�  @�
�9�ڜuF�K�ӆ��K��:`�+�Wv�d�+�D�vw��*����@���Sݿ{Z�zj� 0*3���u���������_�C    hvѭ=s�Y!�?s.�ĺ�h�+�[+9� ��ҹq��}ٍ�����;�?�Agc�+bݦm����;�ݚ�12`��6S�����5�`� 05�r�:@�Qu��t^WLܜ��u    `�ϼ��r�=
�����LN>��:  ��VF���b�����7�[йpǲ=��SÿI�Z����l��[����ҙ���'{g"'��Št� En� � ��9��m���[�Z�     ��9W��wJz�VY� ����2=�   &bh(�OXgt�(������;й��������ѩ�[�N�Nig�I�:��n�`�g+zxbV̶ $)��� �c���::]Y��X�     ������]�;?��V�8d�t�(�[��Kb  ��w�+Ņ(wnq,�e�t&�x���m�vq�.��hw���iݚ^���=�%힜��  4�X+)T�O�Ԣ�S�ks}�z�����=    ��w��=39������:�����p�  �L1�+�
��!j�)���[/��u
:�X6ï�~|��ߓ��h˨�'���>�D����*�r� �Ͼ+ފ��u
������D����R�    ��������M1���1�9@��!�L�u  ���T�ҚuF��Q&-={��c[*V#�X���k��^`����t��C��x�����;���� �[T:_�B�:@�r���d|��/K.Z�     �@>�G�ͽ*�x�N��ږK�����  @'���By�:�sD��­���:��',��s�}�b�κ��>2�����!��=Ӛ+3� ��P�U�q����W�2����;�c     �k���/�
p.�ĺhG.�+߳�:  �@T:7!E.^)Az��إ�Zw�s0��%7���޹���ƺ����:��A���4DݿkZ�*�� ���iM�T�� �T\���+l��{�5    ��1���s��{�+$%�=@;�CrI�u  ���y��uF爮��~�p[�[�)��cɍ���o]Թ���9�Æ����?�z#���Ӫ��) �f�����H��\��}1Q�c��g�    h]���OIS] ;��|FI��/�  :IJ��%E뒎���ܯN��i��?�p��F6^s�sn̺��2ԧ��^���Z#��]S��^ <V(O+6�� �E��s�Ki�%S����    ���s�8&6*�Q�w���������   Xq�2�X/Ygt�({ql���d��X2������K�S�ӭ[�YOWF����8(�z��wO��p; ���zY��ak������2F}�8�غ    оF^~ٱ!M��69��u��|�\��  t�
��'D���[w��1"�%3z(��������͋	,^����]S���: �lB�t� ��#������/�F�����Ժ    �9V�}�ӳi���Z��c��$�Q�7,�@  @�IK�RZ���,�5�w/ߙ��u
�O6X�6^urt�w$6+,���9:�o��V�6���i5n <N�ك�:��s%���!��ll    XZ��}���݁�s]���|�  :KlTʓ�'J?	��ԩ�S�-hO�����~���oH���)�,��:��!y���3_����JC�N 4�P�S��Yg XY��\V]���p�:    ��6rf~}��PNoV9��u8��!���t  ����RhXgt sa,�u���8h#�}�s�*�vwԺUZ��m��5_���]�
��v ��Ŵ�P*Zg X!1j�ym�udz���     4��mt�P���{�{���J���8  �$�VR��Xgt��;
c����@��e�+��3�]��[�Y.������v �~Št� �Ժ���|����3��9�    h�^����^��H���������   X91*���K:Q�ug^0q���X���0���2�q�W��J�v�t�ak���X��1� x*�<��([g XV�,�3��.��9?a]    �b���_�.T�o��=�=@�r�}�r�� @���z�:�C�{2i��{n�u	��X�u��9;��d���W�t�ZN�c�n <�X�(T��3 ,�˒>�d����=�9     ,��3�G%N��8��uД|VIߐ  �"�u�R�:���/�򯵮@��I�r��O�j�燒�n�����Ç��x���R���w1� ؏�*�/�+ڀ��������̅��/��u     �e�YW�J#V�*��HJ�{�f���Y�  :GZ*Ji�:�c���y��-���@{`��2�iۇ�t�uG�;t�_#�s�h1� �@��!��6U�⩝?d�    �J9�cB���Aw��9��!���  @g�sk����]���.A�c�6��uI���n�v֕Mt��Cr|J� �jC��b� �_�6�X��� �T�k(q7�$w��M���u     V֜y��>����
1���J���x  �Q�ܸ��܊������s��;��-hm�: ��%�5b�}�:��p;�Tm��ln �_L��9� K#��_v]��,��od�    ��&wn�Aal�F��s�s�J�K ����   +��e{�#:ZT8e�M}ʺ���Y,�Ȧk79ſ��hw}=Ys�uZ�� &*�/J�n� E�o�Lr~����f�    @��p�
�^`�X��rI�:  `��T���uE��>I^3~�fM�h�〭=����#I�Y����T��80�z���R=�j ���ʌb�d�࠸�F��c�ۭK     hk�̿<F].���[ 3.QҷV\#  :AZ��ҪuFg�~:�t���o�����:|Oe�n_v��,��8`�F�}�n <�ب1��4��䕅���b�    ���ؙ��0��T��1��{ 1U��ZW   ���k� V7b��K�u
Z�8 �_u�I�{�uG'X���:-��ݿkJ��� ���Beں�"D����
�'�R�e�?X�     к\,�����G��ϓ�ǺXi�^RLk�   ��e�%�\���>w���-�hM�=��Ȧk��Y���U�]z����hi��oה�Նu
 ���b�b�`�4)��V�uŃw��     �Ď�pewQ�?��%NqȺX1.QҷVr��  ���s��9�H��t�p�拿a�������k_'�ʺ�{ؠz���hr!Dݿ{Z�u
 ��z���@Kq%�}6����S�5     ��5/��j�����-����\�W�g�u  ��
���q�
H��CQC���9c]���د����`��7I�ߺ�ݭ�����^�4����h��v ���ByJR�.�T�������|쒯T��N��    �*��Q-�{�='��.�aE�$'o�,�P�K�r>c]  �|�WL�RL�K�8��������6�c�F7m�ZҟZwt�c[��n^ ���(�d��) ����RZ�� �Qr;|�9��K    ���}�I��?,ų���hg.Q�7,9�s  ����-�C3pI�k'n����h<��I�����]��&6�/���n��+�?���,�< &����� �#�}ù�=����պ     <��[_]��S8ͺX..��ϭ��   XFQ�ܸ�u$E�I)wJq��[���qO":�)1ܾ"Fs�	hr��n ���9� O&�{��7Ƕ�&��     4�­[�Z˟�}�)�?d�,��(+6�  �3'�e6�Y8�5r�/J���xJ/�	�۸��t�uG'��e�n��:Ml|��=�%� @ˈ
�))��! ~Yt{��Nz}��?�w�     ��J��yW��n��\Q��vR�u��bZ���$ǌ  hS>Q�3{�,��=��f�r���M�47�P�8������K$��N��������:Mjj�����Xg  ZH��*��3 <�/+�*]�'����u     X�5/y�j��]��!{�{���2=�A�  �e���RZ����D���u=��/��u��x��s�����"�NНMt�ӆ�3Ф�+uݿkZ!F� @��iM�T�� �s�����
�\��u     X�g�J|�L1�Fܚ�6�{V�es�   �"��
�P5���\��i�p~ٺ͉w<ƺWm���臒�8��62�����x�Z�{�Tn ���OH1�. )�}�gܟMܜg�      mjhC�y�����_�n������  �e�ΎK
�!�E�����f���Ā;ct�5/�WXwt�l�u��r|
�Kꍠ{�T��/T ��ӊ6��F��ű���%     `e��������?w��b��U�7$FI  @;
�i�:ߩ7��|��;>��:��[�y�{��/f�}��2܎�IC�{�n ,HlTn�G��
�'��p;     �e��K�\�w'D��\ѺX�PW��YW   ,��Y'��\L˟[����Z���0^�}^�ό������S:A�N8bX��#���Qz`��f�5� @+�A���9���F篕��8����     �ֽ4?�H�a)�^Rb�,���e��3   �\:7.��:����Ή�ϲ�@sa���u�n{W���uG�X�:�Æ��3�d~2>��يu �Ť�I)�Zg )Fw���:��»�[     @sYsV��.��t.�ĺX0�(����.  XR�:�X�ƚf�3=o����Zw�y0������Y��!�Nq��k���Xg���,i��u ���ZI���h`����һ�c�ۭK     @s[{f��1ƏK�8�`!\�G>7h�  ��B�t~ܺO��ٴ����/x�:́�P=�\!��WL.�p;cz��p; `�bh(Tg�3�N3��+��x��     �@L���Rػ�Q��(W��TlT�e�  ���)鲮��a��k)EwC�;�ȫ�=݅�o��Nq�U���@�(U���)��S  -%*�/J�nt�U���e�˽w����u     hMg��v5�9����)k�<5/�7$�Y�  �G��*��x�g�9�㒫�;`�����k�.�7�K:E&�:�a9>y�To����`� h1�:�X��� :��)Qr�ޱK�.     �a���)i]����[���J���x	  h1*����Vs��Iw�{o|��v8�@:�Ȧk79ſ���$���:d��:M ���vM�Te�. `abZW(�3��眿Oޝ7q˖��[     @{Z�a��Q�����[��q]�����   K&��e�<��V�����s
��%��q��/u�\�+���[:��F�I�u��O�g5[�Yg  ZM�
�I)�,?#��<�?K_����k     @�*����˧��޺/K�y�����'���.9ψ	  h�3���b8�ow�|�����)���5�i����a�N���KO_��:M`�dI�'�3  -(Tf�%��]Ey��ȾsⶋvY�     ��2x��L\�c
�U�{|4#�(���  @;�J�&��Z���8_Vw�Y�x?K�:�h��+G���#�i����������nj�����Xg  ZPlT�mo�����˼c|��_�n     �m茭/s.~Z
ϰn~������3   ��Z��|��{�su�&N"t ��v��2�����I�r�w�R����  ��*��Z���K.�x�Ng�     4��[n+�}��(^����~QlTk� ���9�<��x�P�ދ�3`���s�9!����2�-�d���΀�FtϣS��9L X�P�RlT�3�v�:�>_w=��qW#     ���~��#W�<��&I�u�����K��!   -���B�:���%���6Ϻ+��3�iۘ�3�;:ͱ��Qo7g
:���5S�Yg  ZP��*��@ۈ������7�k�     p �6�礫��,�@��%}Ò��%   %T�ks�x*>���a�N��o�[�`���AF7]�21ܾ⺳	��nWq��v ��T�2k]��(��K��o��:��     �������\=G.��(W��S�ʌu  �As����8i����Yg`e���S�0��w9�d��i���`�u�L�W��^�  '-��CR�A��!�s�҅7}�#     ����p�H=�>.��YhS�{@���:  ࠤ�)���E�p=ϛ��=߱N��`��C�n��O��6�Nt�ӆԝM�3`�RKuJC�N ��P�W�2���_]&����     ���q��%w�s:պ�����%Y�  �E���2w_w��+': S�`�9�p��W$�o��i�z�lo�g��    IDAT�P!Dݿ{Z�F�N ����+��@ˊrS���8��-��_�˺     `�������׾���G��(���z��Йb�&��I���  �59�(�K�8 a$7�H�w�k�%X~\Y�|O�bɭ���Dkx�ԩ~:>�J�a� hIQ�2#�@��sA�9��g��$     о��0�s�vɝ,�,^*�BL��Y�  Z�O$ύ4-#T/\�{�8�:ˏ#�mn�ƫ�]r�8��✓N:r��ǬӌO��ha�: ТBe����"��]�ɱ�ߴn     �0r�egD�W���nA�q��]}�   �j��Y�(��V������,6����2��&�{�n�@�vn ,Nl�n���%N�U��    @'�yɭ}:Q.�Pr�hĊ��Y�F�:  `Q|�˖��Y��wYg`y1}��F6^s�s�;� ���G4<�|�$Q?~��z��a �E�A�|A��u	�B�-J�\���G�K      ����<2q��)��a݂�%}ÒcD  ��t� ��uXR�I���[�w�u	�Om��L��ͬ�uY'`��t|��v �����������(����ֳn     x���?Tؑ��}�):�����*-O[W   ,�˲̶���kۭ+�|~nS#�9C.�غ�S��d�����$��eM�W�3  -*�ˊ��u���kH����;�8���:     �ٍ��rCR������{�,���P���   X0��N�B�ڋ���o����p�X������t�uJ�:t�_#�s�X!�j]�>:��K  -)���:�� ���k��������K      Z����ω>nw��Y����ܐ\�[� @kI�R�[g`��SI��	�7��n�,-VL����F_�p��U�<�w�4D=�w��v ����i1��G���%�*�m~>��      �W�-���sݳ��y��{��BeJ
�u  ���Ž��cij�u����Qo�|O�T���#�[:U�;��[c�����M�W�3  -*�����@s�x��2�3�i{     �%����.�6�Y�-hc>��wXr��  ��CCa~�:��z^=����u	�Omft����#��l��>�[�k��0>]֣�9� @���`\��5 �/��O���O�m�ٺ     �����uc⧝�!�-hO.�#���   8`����X(����������u
�������O����n���:+�TmhW��v �bE��n~It�̕����3�     ���wl��gKϐ�ՒR���ب(T�^  ���N�b�t��\��:K��mdtӶ�Jz�uG'�&^'9l��eB�=�N�R� `qBuV�6o�4�m��G�c�}Ϻ     �m�?��p��N�nA��A��  @K�i]�T�����$��ޛ�w�u�m�Ѝۏh��ǒx"4�f�GG�Xg`�=R���t�: ТbZS(q#�s~&����s땒�Z      K�]Cs����>��w�XB^�oH�g�C   �R:?!���"����'�;�Ϊu����h��b���@��:�l�\c� �x1*���+����#�:����O3�     �n�׊c�-N�Ӣ�7�s�N�ByJ��:  �)q�L늡~�df��<6�����l;E��',�;��ae~�*Q?~��z��. ��	�i�:��(7᝿xb���-      x2ѭ=��?
!�s�ںm"�RһF��  �fӺB�`��E��ה�������к��$npi�B�,��vgnos��2� X�ب2�HrQ7t��D��     ���;�l������A�Hk
��
  ��rIVr�u����Ci�uGb[���k~�9����֭���5}�X&�ي~:>k� hU1(����Ut�������-[��:      7�!����	'[������.�_  �+Tf�%���������Zw`qX7��s�n�>�.�,�Z#��u �������dQ�!4r�1�     к
c���g��r��-h}�:�بZg   <)��N�AJk�O��x�u��-ld�ug:����tґk��D���vMi�\��  ��X/+T��3 Q���Ͼun�n     ��ސ���x�S<Ժ�������u  ��Jg�%�̮�ez��p�o���±��eE�b`{{���u1�ަƧ�� /�
�Y�
�B*��z�W��p;     @�)��oL����JrL�`��Bi�P @�rr�.��F�uk_�߶���1�ۢ֝{�c�c݁}����u�X���b�N ����4)�5�`�����a���b]     ��7�!�;�q�\<ƺ-*�RһF��  �fÍ�m�e\8|�d]�V6ݶ6����31ƭ�����LkG��2� X�P+1܎��j���>z*��      ��0��߹�էH�jI�uZPZS(38  ���t['`)��3����u��-hݦk�宷��>�9=�r|��Ja����g�3  -*�u�RQ��1~���X�-�-�      �93�[!�ϲ��Ჽ�=��3   #�/H���-�'e��2~���Z������������K�;�s�=���L���0g� hYQ�2#����kH��B�?��v      ����g�ܯ�ܱ@�^R��[g   <[��DHs1V�[g��1��bF7n;_N���ϭ_ӧukz�3���3����u �E�ʌb�d�,����8>v���[      �|�n���cL?�6w,�����Xg   H����XN.���������%xjlpo!#�����;�X}=Y�,��l��v ���F��v���mm/�g3�     �'31��kls�b�ʴb�f�   IrIVr�ڶ�(��O�{�G��K���Ե��I���9���u�H���ȕw �E�A�2m],3�#e�
c�w�<�0     `����ra,�N���(�{�{�*�BeJ14�C   $I.�m��%C���L����Sc��E���k%w�u+ו���:K���i��  ��P��"K�Ц~���Я�
��e�     ��2�3�u��cAbP(MJ��o �=�0��Vj�?~�ǎ�����z�E4��$�ʺ����G�]̕뚚�Zg  ZT��e�`Y���c�M�^�]�      ���o8�,�k7\������c����b��4��wh���   F�mpw��u
��S��Z�JI/�n��c�{X���H�m�x�\w�:K F��Y� @�
���@��r�����~m�6��     �4&�6-7��9��控�J�Sb�  �rNJ�l'�Q������+�;��poI��I9�<^����`�TI�:��  ��V�%qE*ڍ�۹䷊;��;�׭k      �^���rag��N�����A�K�
��
  ���mqG��J�O����X���1���־r�!Q�-�x��;�t%�8H�F�ީ�u �E�ڼ�֬3�%�s�3ewja����     @{����������Xэ����Bu�:  t0��Ph9W�{�u������n��)�ͺ�ן���C�3p��=���� ���i]�T߹�]D%?��wn�'�      t��g�ω!n��z�4/߳Z.���   *��bj����J�o��=7�����ܛء�!�?����ue�p���� )*Tf�p;�D��_��3n     ��������}婢'*3���  6\��:K-�=iy���x<ܛXçI�^�&���Z'� ��H�+�  �*�R�[g K���$���3���X~ƺ      �mz������I�Q���A3�
�)Ŕw�  `幄q�v���k_�[w�poR����#�F�<��n6�����%��: Ђb��X/Yg K�ݒI���[.��u	      ��
c��rI��Q���ByR14�C  @�a�{��R�z�1��Ca��I���,��T❺��u���*[g  ZQ
�i�
� ���
c[��s{~�u      �D
�\�Hq,�R�?�4o݃&�BiR
�u	  �$�K�Ÿ�(���OgJ����1�ބF��~t�{�u�\O�I��]�9��3  -(Tf���r�2���eN����%      ���عe���N����nA�������  �����]��z���Of݁}poF1�,�	�&����U��55W��  ��X/+6*��"�r�?�0��ES;/~Ⱥ      X��.���\� :�5�լ{�DBCiiRb�  X!.À{ۊi�+W>n��}�u k�U��p�poj��kdu�:�p�S��ԭ3  �&�J�����������7_�C�      �`�l��� �EI'X���$]Jrk$�  Xf1(��k]���|�����+��W�N��&�2!/�ۛ^O�[��\��v �"D��i1܎�J��!7���     �.��.�^��Y��Jr���>iMiyJ�� �2s^�Y�
,�\�6�99i�@Y���?��	G�+Ï����_Uo�� �0�:�X��� $:����Tܹ埬[      ��v�ֳc�����-h.��ϭ��   m�9�v��2}0q���ƺ��1��DR.?���x�p{�.3� X���y(E�q�})��L��     ��&ƶ��;5*�ͺ�!6�
��  ��\�e��ec���l��ۺ��%��g�Uۏ�>n[��^�+��U=�X�4D=�wF���  �ByR��B˘�1�Ӊ[�V��b      ���=wΕ��}���nI�#)k�c�.Ir�  ��p�+�J�XN1��eU-����[�t*�P7�$I/?����Ź�V�w��40� X�P��B�:8 Q��i���ߺ��-      ����[�;�N�ܷ�[`/��j��  �]9'%��lw�Q����k�[wt*����ۏ��j���,���.[g  ZLlT������jQ���s�[S����      ,M���]ػ�ף����&.Vgy�  ��K�-���F_�L_n�ѩ�u �u��}.Jo����9r�*�u[g� =R�c� �0!UZ*H1X� ���=J���m�oY�       �f���o�Q���n�-����Xg  �6ӺB�`����4����x�X�t6�[��G��8p]6���Z#�0�p; `!���4��hv1�_��[u*��      �ߙ�z��i�%7X��V(O+�5�  �f\�#� �I�W?e�щ�t�.s���u\w��V�{r^1ZW  ZI��K��F�r�蒍ű�[��|N�      �1uc~jb�Mr����u�D�ҔbZ�  m�II�:+ ���}��ϱ��4�z�5O���;p��xg��P�����Xg  ZHLk��9��IE�o�_��=Jһ�����Tu�=�If&٨���o��!@4�8	!r[n��LWѳ�+��@�U�(A&�=D����芈@��LwU������}���	�LwW��.��99�9��;��Lwէ����ק��ػ      &���/������-�Z�Tx�  �J��	�&���W��1�M���Q9eo���pCd���Ccv���v ������xV�����=c�p�.�      `���bm�ާY��.)z���%�f��;  �Pb�<.�螹����zw�NQ;9������I[�[p�v�آǞv�wE�H��Wk� ',�dO���1�;�M\U?r��x�       �b��מ�,�����n��PR�}�BV�.  �Β�ʬw6K61'v~�a�;ep��I9�7�q�Й,�%3�� X�[��1��-y��D��      @o��L͔&'Д��wXTj�K�C�  `�B&e\q)�SN�k�3����NS̿$i�w��Swj��m�xEL����J,� '�R�ԨKJ�)�7j�~�:3�[�!      ���{���6�;d�7��M(���)+y�  �!��K��靁���c�����ڻ�SF�=��ĸ}(q�}��-�� N�)�Ÿ��,|Z�ē�      ��:=uS&=M>�݂MfQ�Y�;  ؐP��X�bk�i^�1X�n��ܰO
?�݁��`�>�b2ՖZ� �!���Rʽ3��B�tc}WxR�����      ���t�����'*�~߻�̢bk^2��  �ub�>~��U�_�k��1����&���A��݁�)�x4� �-��� �Ί���0J�ߪG�;�      ��c���!�ŧ^xݭ��
i�w6I*��*m�#�� ��	Yy�{>07>,��n�m�.�Ne|g���^�ۻ2�g�;�~%�d��T�z; �DXRj/zW �$��7��      ��v������K��[��R���;  X�P��N�&��{������Q�Zwe[�?m���O��)�
<��fGy�� �G[��@�A-do��Ω�T���      �u��~�6{��,do�/(�F�  `�J��tI�Yy�w�(c��I�<��-K��_�t�w�g�DI���N������Zi�� ���Yg�;c/�'�~�vt��%       ��*�Mf����-�$�I����  ����+5k��tA��ݗ�~�u�]2���I�v�_&��Cm�̗ˠju�� �Ge1�uV�30�����1��v      `8T�+�$O�e�݂M���y�̻  �P*�{��ȔR�m:�R�.E,v7Á�$��;S.��2���-� �����Z�ċ�p-do��~�ح�Y�       'n�h��ڮ�=�B�v)$�lF�  `M���qGVt�ܻ{�˽;F��x�-��;�1{woӷ���;��_�)�� ��ւ�h{g`L��=Y��d���'�[       l̾�?/Y�{��y�`�����d1�  �&�e9�Z�Q(M�7��=�_��n%���;&�w�
l\9��e՗ی� �(u���Ɣݚ��1n      F�����!m�!)��l��Ql�X  ��B6� '���l��;F1�Ӯx�s��w6�Swj��m�x��}��N�3  �bW�9/^x�f3���tp~��ۼ[       ����Nm|�Wd���J�9�Pުl�n1�  �b�Ԭyg�K�X,N>�;?�y�Q�I�>3�7y7�7��T�r�˸ ��,)�Ÿ���.����      ����X����Y�BY���AY��;  xD!+�Í1�w�W����>�w�;�!�l��F�����.��  ,�%�P�lᖴ%���t�/�K       �_���ǂM>���w�,v� ������+�)v�+o��1*��QP������ɣ�[]� ��J�)v�30^�)��6S�h�Õ�       ����_��>Sy�)�N
ɻ}��  <�Pb�>�R��Ӛ��;cT0p��W��$��wz���`�]h�x�  �,ve����p_�Jϩ�T���w(      �X
V��Le�|�)T�k�G��؜oX �o�wt����������Ĕ�,�E��_.�"/�V�� x��Z��'f�����G�>�      �������\~��ɻ}��-F�  ��Bi�;ެت��A�Q�b�N;p�w�e��-.���RK�
  ��[�E����kg��=��_9�      `p,>����gIٍ�xcsT1r  2�_���o<ƻc�1p���K�Y#&c�>b2ՖZ� ��:+R�zg`�4����L�jU*ɻ      � ��o浙��!�^(�%��	#w  ��B�2��cϊ-Y�5�1���طx�)�^�݁�c�>f���  dEG�mxg`,d�`����#��z�       |�#�?4��J�w��I�*6�q  H��;$)�x��7|�w�0c��c]uV���^Lܽ�ERu��� �IQ���]��g!���v���+wy�       ���g��<�	
���[�')Wl�3r  RV�.�@���a�b�����mm6[_�t�wz)�    IDATs�w�ػ����w �72�F]J�wF���J?];r�7�       l���}����
��݂>�&TھG
ܛ `\Y��HV�rԶ=�_����w�0�;�j��/�����v�"��̸ �@��̸}�}&d[���      @/T��n�D��p�w��K�   +{`PXQ
ݕ�3��^�T2�^�<��ݽ��yW  ��-Y����(�?.�gU����       ��v��?X���0�݂>`� �XY�;�b������zw#�=���N{�L�ٻ��w_�v��F�; 0@,�J�%��(S�Z(��6=��n}Cû      ������3��J��J��=�1F�  ���I���,f����:0p�����	,�ݘIwWW�3  �ĒRkA��@?��2�~�>=��       �.Xmf�R��BS�zנ�R�ج3r `���:�݋N;p�xw��z`߁��t)<ջEե����; 00����٠B�wab��3���;      ���=�KK�d
�ϻ=�
F�  ����]�Ab1��!�a���B\oqf\��PĤم�w `�����r��Y�jM�S��/��      `�,��yR+<U!{�wz,����8� ����;��\�����w�0�h��x����ߐ�[�_����0v�:��f��� �U�ېu�=��+j�So՝�qB      ���;o+Z����[���ǂ�GT�nB����(��(nQ 0�,�R�x��e�����O��wɰ���Bx��uyp�|���� ����+�,{g`Ԙ�H��Z���}�       ���t�=�P�QS����ĢR�.c� ���mx�w�8������1,�*ڀ�ܰO�yw`s���}�1�k�� ���T(��30bL٭Eiۓ积�W�       x�ٙC=�����nAYRj�3r `���X.:�k�+��Ha�5��zw`s0o�<���c��  KJ�yI����������y�G�<�       �ح�����=�B�v)�B��8�އ]�  �/��;���O�r����1��ә�߰E���������Xht4����  Sl-H�C0"L�j�.��T���7w       �͗��t�!�^$<{d��^t�C  @?0p����̊�/yw�봸�t��ӽ;�y����n�t�ܲw `@����^�����*�U����       kU�>��Hg���-�Sj-�r� 0z����Y��l�7�'�A�W�:�^�݀�UD���Of�]�K�\� HJ�Y�������4k�ٙ�_�.      ������R�����-�Sj/�  ���x$VlQ��F�AǗ�:�v��ϲ`��������N��;�xg��{��.4�3  ��R{�;�!����g*S�!       �;N9��J�]#�GDزK���  ��JͺwY6ќؾ����|��wʠ��uH�~޻�//���/K�.�v �$Ɋ�v�),�L�g�      `���T��R�
I��5��,+uV�3   �R�=�6^�1���Ѿ���t�w6_���	#�ݍ�kv�; 0 ,�J���������G�;�       �2w���rv�)��wzú+J>�  ���E�=n��1���Q(�׊_����2p�"&}�آb2� �3K�Rk^&`�,�H��Y�3��       �V=\����ؤ?�nAoX����H  Í�N@�w�;�?�1�����|�;N����UI;�[��&J���zg�3�K�-h��{�  �Y*����a2lH4eo��T��C       `�Y8�k�G����d$��6e�N�8 >Vt��Y�&�;�}����/k{�.����ĖW�q���cR^$��
�v ��"�vl���J�0n      0��է+oTVz����k�qV��Z��,  È?�qb,�{��՗xw"�'��JYA?�_+mٽp�|C�%^S��gI�Yg܎���,������a�       �V;2��a�W�[�qV����H  Ã?��)uߠJ�=���r���?�RI���V�;a��-�tl�� �Ƹ=`!;&[O�N���-       0(����D̞h��ڻ=;��y�x�<  C��;����w���΋�;��~޻���oHm��{j+�  o���R*�K0�L!{[}z�yՏ�m�;       ͱ[+���{�)���nA���{+�� 
Ɵ�XSjw~ѻb��a���w��̲Oyw`0�y��ڱu�;c�,4:�kv������q{�]�����e��9�~�       �\p�Jz{��aJʶ�Q���%  ����,ozg`�d�v��]�W�%���' ��j���r�;a�ԗی� ����>��ٌ�      ��է���&�3��w6ȢR�.��� �@�;�,�:�7{W��+o�+�
���FG1��>Qs�-}un�q; �;��ذ�S*M<�~���z�       ������d�IR��l�%�漬�z�  ��a)z'`Y�w�e��>�A���Q�_%i�wGL��b�;c(�o�ڊw ��%�f�q;�/dأSή�r�׼S       `X-��i���Q�lTRj��r�@ �@2�X�!/��;cPv�����z���z�`�����}̩*e|	=3������0 c/E�ּ�
��h��Z��Ly�       ��p���V��A�za�.e�;�3  ���W�yW`HYV�f��|G���o\p�C�b1n�C��tl��1��"��.0n ��ۛu��X+Yi���      �ׂ�g*S*e/U�x|���βR�'� 0(��6 �bR���;�G`���n���[li��{g�F;��_�W�ͯ �����<v��E�)s���w       ���-�߳�=[
�y�`c����^��   G �a���{�o�������a�~�=�ҹ�lw�-)&��ե��x��S  �,�۱�_�){r}��Y�       u����6������{�`c,o*�$�a  ��%�ؠ���R�����?���I
�ly�t�E�1�1�+ǖ���l|  �Y*���۱>!{Om�㞽��J�;       �E�c�r�]���t�w6Ɗ�bs^�y �#.����ϪR�7�p���8yrr�ݒvx�`8��}R�=m�}E-4:�ZuEW� �,�J�y��sk-��T?R���!       0�N���7��/K6�c���M��}��� �f�+sD�w��؇^��/|'��LN�L�۱Kͮ�2�46��W/�/�+ǖ� $1n�X����<��       �6=�����X!ky�`R�بɸ  ��J�q;z�;��yWxb��M,��OyW`�,6:���u���*%��bK�����F�; 0 ,v���۱v&ݕ�윹���       ���-S�R�#��^�l�E��,��%  ���E/Y̟���;��ᅁ������%}�w�S�[����k~e���fR}����]�=��1�T xtV��q;�*�c)dO��>���%       ��>�V�Y2��0���{׻ ��`��;zȒR����^�?H�����Lw�.�{����}�k���ܲ��" ��h+��%��'�Q�>P�Ξ����       xh�+w�������-؈�:r/��!  �<+�Pz�ȯ��K�y�w���w� 9��M�I�n��@^$՗��I�&���U�j�m�5���R[Ed� x ��J�E1n����֧+?����c        ������n���}�_n���{�~��Cyҹ �eI�Y����I��l~���]�نgq�	�,�J���c��m���y�qς�W:��6;��[ֿ�U�=�usvg �o�:n_�v�M�
�tU}��F�       �Z�OWި��3fʽk�~�]Qj/��x  �=���oR��z�M���1��έ�w���$��N�hʋ��FGե�Z�B�L�R�R\���Bե��V]��BK�n��� ����Yg�;��¬�tAmfj�;       �>��?���|��X���ݻ�r)E��)��  %�7�Txg`Yܹ��}��[?흲��N��}W��@0}л�gۖ��o���ɒ�o)k�DYY�F�fR�[����h�Zi�*b���/ ��I�Yw�;C'�lQ.=w���/{�        6n�y����E���n��&U�v�2�  FB\���-�#�&��z�5����L܏���W�g{w ��e���rI�r��R�r)�dy�?C
A�BP���L1��UĤ"&�ER;/�ɣ:ݨd�g �]j/��w�N�eK9\q��
��       �����މ��4Ȟ�݂%e��(de�  ��ŮR�����s��fo����.�,�%��ߝY�9��  � ��Z�-��k3׾V
|�       Fс���O�^蝂��m'+�&�K  Z�f���~�����Iʔ�Z��  �L����k-�__���j��       0�n�tkӕ�Jo�B���:YRj���w	  C�
�E��ؽ�K޽߻c������/}�V�^��  0P,)����.�P	Me�ק��w	       `sԦ�~U^",���)�d].� �VVt%�~�`�DJK����,c?po���K:ջ  ``XRl�K��]��rL)<�v���x�        6W�h��!��3��݂�K�%���w  C��w�H��W�R���X�M>�^�   00RTlԤ�{�`�X�\����*�       �Q�9�Y��4I_�n��Y�Tj-H2�  �%Y�Cl��b񘽟�q�w�f���+���
z�w  � ��+6�E���Tl;k�h�N�       ����[�0��O����n��Y�^}گ%�  Z�[�Ca�\&���zWl���+駼   �]��<�v�M(�~�����M��)       ��p��[�v��L)�c�l@�FJ�w �ñ����|��~�;���o%� /���A�w%m�n  �dyK��(>U�5�Jv�v������8�       x��;o+Zw|��m��W'�S�{�N�dE[�4����� ��dEW�7�30�,KY�m}���.駱���e��N��   ���X����JW�>v��x�        Y������k̔{�`�,)5�eEǻ �������'��ez�M��4�w3�ܻ  �Sj/�:��.s��t?�       ���ԻK��|)[�n�z%�ּRg�; ��`��"��K�}{g�»���r�~���~Igyw   �0�ւ,oz�`����r����k��;       0\�f�f2�sM����uW��K��� �qg��c 䝟�N觱�'��   .,)6�eEۻC%�S�<qα#o��w	       `8��\�ϊgI�3�-X?˛��yɒw
  >Rds��`��}�%�����2v�3ϿaK0�I�  �M��b�.Ůw	�JvxW+�=��_:�]       n�[��j��1���݂�]�f]�
�  6]꬈��` XR�#{�}��˻J�J:ջ  `3Y*V��Ј5!���]|�m>~       艅W��>K�����
�f]�a% ��TȊ�w�u)^q��7l��臲w�f3�^���g  ������Z�ģ"q��B����Ե��N       ��O�f^����'�����%�漲�')Ll� �דּ� <P��Y�,.���^����;��   �źM�ּ��D�B7��ק���n       ��`���7&e?')z�`�L����Y� ��,沂��c ��+��a��)�^�1�{  �+���:K�&�-J�ys�S��N       �����;C�]*��݂��nC�9/�y�  ������R���/~�c�;zm|���V�Az�w  @ߙ)�dyӻC��.M���ʭ�-       ��R=R�hI�7��݂��f]J� ��[Rʽ3��f1˭3rW��f�~ھ�H:û  ��,)6�<k�}>Y8g���O{�        ���̡���֧��[�)_}�*2 �KJ�e�
����U���&|��fI
z�w  @?Y�5>5�51e�謅��;�[        �:��/Lj�YR�G�l�E%2 FD�H��3�G��o���;���Kc1p�������   �bE[�Y��G>�ąP���N=k�Õ�        $龙��e��LS�g�-�Sj-(u�!  ��Ů,ozg '�;�W{W��X�C*�DRٻ  ���Tj-H2���{�Ӈ��͕�w        �h��J}���W���݂���2�c ���R{ɻ8a��sϸ���2�,؋�   zϔڋJ~���t�:}�+����       ��t��6]y�I�{�`c�h+6�%K�)  ���]�R���`�D�U�wG����}���<�,��  ����ب��w	����L�+�3S�        
����Pz�XG��Ul�d1�. �QY�e݆w�fV��{7������ �H��+6jR�@�I#˲K�f*��       �Z�OO�]��2S�z�`,*5벼�] ��3Sj-xW ���=��_�wF/�����/}�VI/��   ��[Jͺd�;C����G�ӕ[�[        X��-��+g�IZ�n�F�R{A��$ɼc  �&���&C,)���]�#=po��K:ٻ  `�L����^/�a-L�n)�H}��w�-        l��_�X(g�J:朂���؜�,y�  �,oɊ�w�!����	遻��Ļ  `�,)6�e�����Vg�g*��.       ���+���&�1˾�݂�]�FM�
�  d�Pj����=uou�|ف���x���xw   l��\�Q�b�;C�,�۸Eg�����       @/��r������쟽[�A�uY��. �33�֢$�,��`yg�����=��%��;   ���Rs^�蝂!c!ݾ�g/|����       @?��2kҹRv�w6*)��:<� �#���{g ����i�w�F���]�^�   �>��YVj/�Oc���ԟ.���׵�K        ��Lei�N9O�>�݂���RkA2�N ���Y�I"=Vl-uxgl�H�O{�;�����   X3K��yY��]��cR魵�k_�J�OF        ��3WwjO�e!��z�`�h+6k�Tx�  ƀmY�'�`D��E�	1�w��%�   ke��بI�띂�-�^_����;       �MW������4e�y��R�ԨsM �Ws�֒w�7�����m��5r��;��I�.��   X��m(5�E�3�e��OO�û        O��ʔ�����N�^Rj-(u�� ��Z���#�RV�+�#7p�ͪϗt�w  �	��؜�u��K0��V�J�V~׻       �AP�>�k�e���»gݕ���w
 `T�)�8@���R����5r�`�  `�X�5)v�S0��%������G�K        $sG�~;d�)4�[�qV��u)1D l�)�楔{� �#���w����X������"�<�  �GcݦR��'��^s!�Ϫ��s�        Qu��o�e����K�b�&+��% ��eJ�E)�g	�IRj�^�]�#5p���&�;   �����:K�x�"���V6�#�#�ʻ       �AV;:��L�\Y��nAXRjՕ:+�% �!�ZK���l�B����V#5p�t�w   �ñx�e��w
�U�nOa��#��;       �a07s�?�,�c�W�[��]Ql�K��S  C"���j`|������i�k52��t�;�]���   %uJͺ�
�)ٿ�=}a�^�       `�ӕ/H��e�s�-��Ql�d1�.	��:    IDAT ��^��M���)��Cw@|d]%i�N� �gI�9/�,K2�)��7���#�n��U        ֡>S��;Α�Oy��G,*5�J݆w	 `@1nV���R���P�>���n   �FV�U)v�S0�,��'�ó�?��E�        ����J5L4�)e�y��WL�YVj-H��c  �q;�u��{�e�9�k1�}/x�K�~�   I��R{�Ұq��~����;o���S        Տ�my�N9�BvĻ�cE[�Y���; 0 R{�q;�`E�B��{H�*�   I�T��x�Jؠ�߮�z�*>%       @�1su���q�
�݂J�R�&�[�%  7��Z��ࡤt�|��q���^�dRx�w  �u�J���r�����t�R0�        F�͗��L兦�7�S�K��^Tj/J��, 0V����q;�P,��N-��#�'j��}v��$}�w  c���J�%I�P�1Yv�6S��;       ���>Sy�I�{���,o)6�R��) ��`i�����.Z(�z7����[Wy7  ��eyK�Q�$�BT�~�v����!        ����u�L�u�豔+6k���� `��x�CM�w	0�,���Jٻ�D����/}�V�]��  Ɛ%�����&�;E��U����)        ���Le*��7����KJ�y�6Ob�Qd1?>n/�S��`�)�O��,�1��f�}����;  �x��j�m��S'+�������w
        �l~���C(�FR�nAoY�Tl�s�
 F�m�f]2���"����'b����  `�p�=��B(������K        �T�>��,�_(Sǻ=�ǏX� ��u�J��t`킊���K��fh�g<���t�w  \mG�eK!Vg�{�        ����>�A�KW�o�KJ�y���E�02���Rg�;Z���}񮳽;����m鹒vzw  ���v�I5%=�zd��-        ���n��S˲�daŻ�gyS�Q���; p�,)6�ey˻z)�^���h�v�̮�n   ����
W��ss���h�c���        �>=�g�ҏ�4�݂>H�R��P ���\�Q�b�;���;�����{�o�ʶv�I���  F��b����`�3髥�mϚ����n        'f���Rv4��z��?By���'Iaho��Ȳ����y� #$�<���}�u��]�p��l[�"1n  �f��YQ�S�����ɲg0n       `�T�\�)��3�p�w�Ê�b�&�=B  ��^Rj/�q;�k��ڗ{W<������  `�X�QlTe�����6�s�V��        k7��lb�9&}ջ}bQ�Y�J0  K�b�.˛�)��
E~�w�#	�ku�U7�T���$m�n  # E�β�h{�`de�͂�=7]�        C��;�������-�lB�m'KYɻ Ǝ���6J�)���,������_{�w�C��n�R1n  fJ��ի���7�g�Q�d�       �h8v��_��tI�{���R�ب�r�G�Mc��^Rj/�q;�R(5��+��܃���  `�Y쮾 �]�D���OOh�Y�n��z�        �ީ�T�Vi�R�y��SRj/(�%�=E �'K�b�.˛�)�XIJ��nx8�;`-v��]{��OҤw  B)*u��؎����S����?��E�        ���W�;��'B��nA�eee[w+�&�K `�nC��@!�"��߲��_Q�Ny����>Y�Kĸ  ��%�βb�ʸ}g!����g3n       `�-�T��l��i��Y*��u�nC0�G,�^m�,��['K�����e����'�  �01�ncu�΋M��}r���~|�ʊw
        ��Õ�B8�L�݂~3YgY�9/K�w 5�[�����)��K1]���P�w���s��!Ί�  �X�Vj/K�S0&���Oj���y[��        0f�^��])�>���n�f
[v*��� �ŒR{IV�:00By��L{u[e�>�74�'��\1n  ��b�ج+��ce����       OՏ�m���y��/�[��~�]��$�DX�VlT��Ɗ�{�l�i��]�.�N �U&YZ�+EY*d1�_�X�!֒d��K�RkA�Y�V�T!�n��|�%��¿x        ����*+�w�t��}»�$v�5Y��.��eiu��ZX�R8)�^���`�;�D�񼛶��$���,�R\��������7�MV�$)d
Yi��L!d�����ߏ��81)*u�_4�%�\A�U���R�p         I:����U�HP�q�l�Pުl�IǷ  I����Yf��0�������FC�����/��C� F���c��ו��a��%)+����A|I!+Ka(~��ϒRg�a;��?�>%\Ÿ        <ؙ�߰�jf�y�`�Lٖ]
ۼK ���B��$E���l�)�����w{�ܯ�pB�]�n����bWVt�>f��T,J1������4~�P(��8��v��}��d��q;        x(w�\�с��OY	J�{�`�XRj/Jy[��'�>� Ɖ�RwE�m�M0LR(�KIz�w�����߰eiW�����- ���b.+��ؕb����)��ʫ�ޏ��!��81)*u�1 �?�=E/f�        չ���t��.�N�f˔m�;��aEg�j��=��M����������0�Ż��3[��^�eEW��U�F�Ri��;���B�m�����v        �F�VʧnMT�%�)pP�Ti�n��]���K���]`#B�q���=��n���"I�w��)�Ի��2Y�Vj-(��*�������LJ�,o)u���5��Y�Fm�˼%��:s�ւR���v�P~?�v        �f�U�Z;�\��;bw�=�nC��	`�X���Re���;��w��q���h๕�;K�v� �Ê���8�ɿ��
��ciu�^tVG�ݦ,v���ٻ�8I�����s���꽧g�F�4ha&`�5��1X2��%�^/�A�B�˵lc_0\r�k�Z�I,1�#;�/c�q�H,�@ �4�]�{-O=�������MU������j��=�|�ݵ�|�_�%39�$7��@a���ٹ}�kܾ1@�Ǫs~\w���u        '�;Bc���:66�,9�(v��Iy*�R��(�4w C���B�Xl&�l�����C�	����>I;b� 0 �6���Wh,n<9b�n�l��n��K���7��K
�5Y�JƓQ�����P����X��x�`��Oչ�[%�!        x���vu����?����B���\���ar��B�*�v�4 ��앱#5�w�{m� Ⲑ)4W:e�֊dy�H[�岬)K�5�kG:o��\���R�g�S���xs���8&���܁��        ������%op�[bGA<��_UY֌ N��BkM����݈�@��������cH^p7sW��  ˚��5��Y�.���B�����벼-�r'fcZ;�q8s�Gjs�wPn        ]u�u�����7ǎ��,��{{cI� 0 k��>/K�D7������CHR;���}��>S��R� ���M��R��ʴ�!`���y*k7di]��S�M�yɹ�!1 ,d�t]��ܙD�m����U�;        ؤ���o~�'��I���qQȎMCvI�c00,K��)�[�s���>���cbx\.��� �e-�֚ڱ���X�잧?�uI�ExR�KJrIA/ȷ��w�!�i�4�	1���U���9        �&W�����_&�7ǎ��L��)o7�G&䊣���,d��Zgx!�-�BxY���cx<&�&v �gYK�zU��H�}��\�5e�U�zU�����Bkuc�w���f�y7�ƒ�y��2�v����*        lΪ��Er;	��
�e���,d�� �j,(4W֫�ہ���=�����c�Ȃ��7�?�%}O� zǲ�Sr�ؾmLyO�7
�G:%�Ʋ,���x[�!d&ˎ/�/m���g�!�
��¡��c�         [�-��Չ��A�;
D�*�W�+��{f
�5�k�v]t= �к"z�����h@�8E!Wh,)4jLt��,�e����S�7^�[������#'�7����!���zYx��x�        ����jCo�����d���t]Nt��B��|}^�����c�}y�.v�ǲ����kb� �M���e�u�dO����\R����y_�j˱�ɲ�,kq�
6��Y�L?�J�(        ��*��e��\���Q0`\"?2!W����3Y��<cy�0 R�Vm�6�Q�6�v�
�g\���ԕ$����;,KZ+S��u�X��%E�o����=�/�B{�ʲ�6�t�K�x�2{�v        00���f��g����` ���Ȥ\�;	��c�vS��F�����K����{��n�mۍ\.����r�֪,k�N�M+Hy�)_�������^���h)���Lʳ��4O90���ua��7�r�v        08n���k+?0��os
��&�5))u��I1v" C���� NJ���(�e�]-����
麬�.�� "Y���鸇���w�<|�4�oh�dy&m)ow
��m[��OT'/�N�\ǫw        0xn����?x͢j����q0��T�^����	�� �e�p�$Y�_s�k���u݇7v OQȕ7��<��8q.�(�'��DrGO}�t�΂,�Ǌ��g�.��-�\r�V���
��       �@�`�Gj�p�9Qr�r��\i��; I�e��b{;v C+inӶ�{�~�c��*��x�����s xj��Ph�����\�t���+�'�sr�wJ�.�C��)�Ǖ�s��Evn����'�G|���Q^�       ��pƵ�����^;�@2"_�+�b'�w&k7�:�v ]�#�X��=���w!Ʀ���;����BsE�5c'z�6ަ);6����\��Qxw�?�N���D�x����l����ce�����c'�H���q�z�Qn        ��۷�\���T�73�i����y0��B�%��|iL�Xր�@�mf
�,��X� �!/�D�]fW�|
.�5�+L��+�o\z�����ym\?�[*i�,         '��*��/�\F��Kᅱ�`��BsYj�ɕ�䋣��l 6
i]֮���&{I���N>��m�4/)���	0Sh��ڍ�I  xB&�7cӯ��-?ǃ        j;���������];���+����
��a ��SYڐeM1j@o�z��i�Q���s�7|<嶽Z�ہ�`!S^�Qn �?|�q%�v        �,���ms�e���Y0lL�55�k�
��ء �(3YZW�^U��dYC���^��Vz~����n�폝������^�B;v  ���Rh�^�p믯�N        �-+����v��2�;���֪���΀ô.Y��
�c����\���Z����\��"ƾRp7'�ձS x"��ZSh,I�E `����r�U����I         �m�3�Zu��J�{bg���S�֊�#�닲v��;[��u��
���]}- �{I�m]�Mm�>|���s x�7���;	  '���륇?]9;	        @/�\������bg�&�r���GR����,Ȳ�B�IG�@1�j�i�*��i3�}���3 xl����Wy� 
f�J
���        ���C��f^(���;6�Ж�k
�jg�tkU���,v2`� k7K���� 0x���������}��n�+bg �ݬ�P��$�cG �I��7���U?�����        �/˷]����4;6����u�FM����E�t]��ɀ�cA�֕����-k��G 2����3z�}�����c� �H���9*�'O �!`�&I���*ߊ�        �ߪ��r��+D�=gRޒ�V�:�Ʋ�ݠ�<�B��|��|�BkecR;�, C�����ܓ4y��b� �2�ƒ,]� �br*�_5���         �Ń��\�_irK��`�\�5��ޛޱ�Y���
���mb}A�Z�B;v2 xJ�����3z�]�];���7�� ��gr�W�n{ם��         Ķpk��\-i5vlQ����ޏ(4��uY����؜L��
�����7�d�dy�p p�,���cW?��^pw��3 �N^�Iy;
  '�䖼W,��cg        G�n��T|���� � ˚�֪B��|�����Bs�)��1d�d�F�}��:�k�t�)� 6+�������w�����tv� $��
���[C ��ox_z�����;	        ����]��·kej��<�I�-k���:��^Sh�vJ�y[��1P,Ȳ�Bk��	퍍B;�L `�0����~�~n�h.	���? ��M��x� �IR��#����Q         ���������()��x|A�SY�>���r��9M
_z�L��e�-�����N �.��vQ'�K��;��u��(� ����
?z��{>;
        ����;��N�OJ.�����ɲ�,]Sh,mL{?�|�ڙ���˲T2~��Y�e�B���XV���|�pg:{kU�5)��g�su��};h��k��R��]w�:,iG���uYk5v  N�����:���I         ���7�����������%�ߓ�ˑg�">3Y�:M��c�98 N�/�;�_��^�޳eǗw<G�ہ((� �����Sn        8y�C7|`��JY
�;��<=6l��I��|���Q��}D��3)Y�%�7���F��)� ����6w�ݛ�<���VZ��t=v  N��Wjs�ߎ�        `XU�*��}e�~&v���Sp�sY���cS������w� ?hl��r�m�n�r=�� �.��"I�ۏ���%��x{[Sh�����1  89��z�P���1         �]u�������_���L�V�8��7�䑅��;��ƬSX�Й����)�@lf�y����k��=�ڛK�n�&i<���V�˲v#v  N�s�?X8t��b�         �<��^��?t�;	��8/�mߝ�F^�s�{���5��If���q9<|���q�C�b ����ON��/��z�(ܫI�{(��a
�eY֌ ��✿y���o�n�        `qV�W���Q?!���Nl*�Q����y�O<���{��9u��������ٶ����;����݉��w���Wظ��p�=<|�	� ��%��z�����FQ
�y�WFl9�� ��T8T��M��o@         ��J�m��]�ڜ\xy�8 $)t�����S�Q �/����(�m�L���/�Մ�
�v ��1�gj�u�uy�,         ��=s?��M]#�/��  ���-<�/��c�����������/�Մ�,kĎ �I�W.�ktK%��        `����������;cg  ��3ӳ��O�'���_$���}�-$4Wdm�� �!c�+iA�y�J=v        ��b�����&���Y   0�̞vƵ��6}/���K��'���֪�M/ 0\L���ܫVo�,��        ����<�
�����   `�9+���K{�M��A/����VZk�t=v  N��#Iq���\�۱�         lU˷]��D�j3-��  �f�z�E_�O���s���{[EH�e�Z�  �$��br����'v        ��n~�/%*]-9�:   ��ɞ��=�B߇    IDATZp�w��K���V�uYk5v  N�o8�k������I         �1�{�Fο�L��Y   0�Bxv���k��ɾ���[���� ��\�Ľya�         �T=t�ϼӏK�cg  ��qn���9��}-����~�lv��
͕�1  8I.x��U?y��N        �Ƕ0w��K~1v   +Ϯ�ua/w�_����Q��69��
�%I;
  '�����^���c         ����-��_�s   `�x����{���v$�K%M�k?`S�F�=�N ��qɯV���1         pb�s�w��ߏ�   ��,<����������~�lj�7%�c' �$��W���)         pr������q�   ��^�޷����q/`s2S�X�B;	  '��iu��O�N        �������?;	   ��^.߿������I�沔��c  pRL�s�4�f�Y�,         x�n��#]#�/Ď  �Ȝ�{Ƌ��h���K������ْN��^�f�+��;  '�����+���V�,         85�V�r]-s���  ������3{�x_
�!qLoNAH�e�z�  ����
�+ks���Y         ��?]9����&�@�,   ��y=�Wk���nο�� ��eMYk5v  N�|�/�~�߉         ݵt��L�6�r�,   �äg�j��eF�x
,o+4z 2��������Q         ��s7}�%��Ԋ�   �gf�j��������.��>�fcA��$)�N �	3S�9���*;         z�z����>�QIy�,   �3��z�t��{å�F{�����ƒd�� \��ma��m��         �?��Ŝ~>v   ��3;K�VJ�X����酽��lBcE���1  8I�����o�         �ڡǜ���9   �GN�m��i�X��w�����LB�.��c  pRL���s�_��         q�U��s�?��  ��)h��^����w�DY��Z��c  p������\�         �ka��w�ܡ�9   �y�E�X���=�~p�L��r`���)4�b�  �$��T�<�F�Y�$         ����r�]+�;
   z��.�ź=-��\����MÂB}QR�� �f�����?ڎ�         ���*����$���Y   �k�^��ӂ��{^/�6S�X�,� �fr��x�­��;         ��m���_m�cg  @��׋e{Zp�܁'ZkR�Ǝ �	3iQ�p�§��_H        �1-z�7gWI~%v   �s;'_����^��ܝ�����agYS��ǎ ��s��8���m7�;
         ���M_rNo6S;v   �F�.���=+�Ͼ��S2]Ы��ag!Shp�2 `��N���*;         ��¡�'��C���  ���ޝ��5��౅�¥�\����)4�%��A  8aA�_Z8t���        ��2���%���s   ����s��f�
�ץ�Zv��"�} 0L��,����S         `8U�*���b�   @w9�s��f�
�f܁�bi]�nĎ ��3�gչ�&v         �����n��;   ������=+�Kzn����m��j�  �03�w�M�Ar;         ��-���D���?Ď  ������fO
�����˒.����в��X�D? 0,���vz�}wT���         `sx�J=)��4��bg  ���rgH��v��\쨵f�^*�bm �ęF
N��TNLEo*%R)��T𦂗
^*�Οi�/)�Zr�F�G��$�'/���{��̤,HfR;�\�N����u�L;Hypj�R����)R�w�� �t�C��ի���j�$         �\����ó���j��wҶ�y  ��9�R�4Rt*x�b���
NŤ�Q.8�TH���JI�[W.:I��:�.(礒7���V�����?Ƕ�IfA���̔�S��������_���ܔf�V�Ҷ�Ly0�B/�]@|N���:�6�owkɞ�]�?C��������i�`-H�E�hb�N��hQשSfOL�S��n4�'���~����;p%��~�3�G��c�O�Y���ʜZ���;��V����S#uj�N��R< l�·���t_�          ؜j��t玫��z��!9+�� ��ђ�h�i�$��x�}���q~��6:|N�%��	�}jN������:�a�y���mS�mZO�9���iP��c�k�M�4���,P��p�!�����%����$��Ƌ���i�d/�L%�XQ��(��M�O�a���jtt�?�m8Z�7�G���~����=���_������:����z*�gN��z۩�9��N9� 0t����޸p�/��        ��m������Ɵ0���d'� D֙�>1�59�4Y���*{M���JN�#N�E�dOos��/���0^���=}ty�#�TϜV����i���2��Ak-i���
��)�#��t���vk���M�lλ���fF��FL�#��d�4U
�*��KOm��fs�S�����<�ef��\c!(<�� [��z[Zo{���ն�J�S~�  �ɹ�g8;         ���C7���+*���M��  ��xM�M�z͌z͔�fƼ����G�Fz6iR�����i�(i����N�-�bӴ�0�4�VZ��f�r�s9�smփ0 �����zRp7�^���c�h�)�fF�fFL�#A����H�x�;�~:Z�O�D�b�	��h�=���d�<�T��B�_�ȜVS��TZj:-�N�-���w ����v����        ���z{��ۯ��/~,v �j
I�m�^�ƼfǼvN$�);m��KO4i��נ��4]���N�q��{8�Z۩V�Ճ�"�b#�J�TO�d�����x���\����?������^�O�K��m����r��i�l*x����^�{
�}�rt�������G��K��>kG���r�i��Tky���
 ��o����T�         [Pu�n_��,�^; lF��D��mw�1�h�������E�Ĵ�Y��O���Ms�jݴ�4��X�U����@a'&�;���u����'/�
�}���rA�1�}̖M�GM�%���j�s*
�[�Ϗ+��e������z����5�9mz-6��m�S�0���ra        �8n�.����|���R�$v V�5;�hǄ׮�D�'�vOx��b'à*%��&��&�:��;�>��Ҕ�릅u��Z���\���v��)�8�s�����^p��_"=��R`�J����c�Sd�9f�14U�N'&I%I�]�?�}<˴m<�YY�<oK��I+-�j�k�鵰�9ߦ� O���+���;*��Y         ��-�Ż�g�|�������;v t#�D;'��L�g����f�hp�;���4]v�`֩S~/�LZiI��M�ׂ�W�փ��߷0��s��ߏ��C�fҿ���,傴k,�=�]c���M�GF���)˲cy���n��d&��NM�j�k��5�p���8&�$���*w��         ���+�ɇ��4; ��B�ݓ^���6�h���(�=�ܤj]z`%�C���+�փ�,�޷ SV�?8�/~�ݍ�~����朮�����������=�g,h����؈���#���v[!t��-���^Ն��F��;���L����?t��          �������͒����`�s�kf�Sh?s���f�vN8&�c(���+A�=����Z�z+�������ڧ��n�U��"�s^��;7�J��g<h�x��ƃN��*��pI�DI�hdd��uGK�c�Of��3���B��H��p��uϔw [�%J~�r;         U�`��WU��B���Y ��F��N�Jt�L��3�t*rx6�ɒt��wx�-/7��WL�Y���r����,���)3gI�J����\���#+��uq��P�N�V�Lf�3֙�~���;
������n��e�L�R���z����z����a ��z����1         �'3{��~�Y���9 ���J��Nt�t���%:m����ڂI�u�wV�\���J��Z&3���go\������X��ܗ&
�x�����N��;t�dgB{����B��B��r�,I23��m���vO����r��u�ֽ\K��@1 C�9�¡�$UbG         �T�2{��߻����� �S5>�謙�Ξ-����1����vN8�H���:��V.ݿd��R�o/�:��)���I�D���Z��w���GK��i�x��A{'r��O�9�R��R�$�Sx��\��vM����Vm��������z��z�����'����          C�R	��T^����H���q �D�ݓ���^�y��N�trtځ�2�Hlw�`{ARA�FT�K�Z
�9��K��mI�`��խ��Zp���{����\gN�:s2hz�p*�sǦ����J��,�d��S�.NS�����zp��;k�Zw�T�����;*��A         ����m�����5r���� ��y�u�T�sg:oG�Sh�
�d��v�K;ǽ���K*��(�Šo-�1�Z3��x\��Z��w����蟉�錉���r�3�Sh��
�Si�3fR=�������}k�龕D�m����L�r����*��          OEm���WV��_K��� &G�=��ق��HT.��mvT��z����RC�����L��r�2Ὧ��-�;�Îzg�h:{�3����\3ent@lG�ccc23�i����ΚI�¬�Z��۫N��$:\�<T�;3���ks         8�*�8{��~�Y�ǒ��y l-�{�Nt�lA�v�s��$0hfF��Q�g�)�3�}T_���f-��˹-&���3�޵����$��Cw9��n�����w"�9ӝ)�ǂ����!(MS�Z-�ig���뉾�����Di;!���\�C~'v         �[���=��;��o��uֶ��ߑ��]��;R@�-6�{�����V��<P��&᫵O���n��ź��]�}x]�h���zfʦ�3]�-�ɠ�q�����,S��R��R;�u��u���}ˉVR�^����s����         ���+�Q
o����39���ق�����{%�z�M)��+N�.����L��B�X���|����V��w�x�����^�@��$��s�3��1�}�H�،�s*�*����P��j�tֶT��S-4��[�o%�R�g� N�������b'         ��:��Ϯ��cg0�v�w
��L�k�ǎ�
^:w�t�LARAk�ӽ�\�Vs�W��J۱#!�Mz^A��)�֢�q퇾�;�ѭ�6��A��:g:���\�.+������Z���4U�!ݿ��+^G�<a�T��LzQm��;	         �+�W�k[!�>/i_�, �϶��.�U�3v�s�����I_��to5��j���'�Y{`������ӵ	����2���Hb:g:輙\�M�gJ;��x�U.�U.�ef�JS�6�ҳ[--6�o,'��r�E&�81�骥�)�        `s[>�k���+����uNӱ� |�&�z�΂�������i *��&��&z�y��e�S�{!ӷ3��Lw<��������-�ӝ��}�Lٴo[��3�J�8�9���hdd�X�}�LK�KS��ҽˉ�]J���N
` �k&.����7�;
         ����]��������rֵ.��c�X��v���=�����q �ɒ��Ӝ.=��<���1}m>�����$��G%���tq�{�k[|���Ѡ�fs�?�k�X���� ����Sm�����Z��M�,%�{��F;)�a��w9t��b         �����|jە7��7�^�, �x)Ѿ�]����g(���K�m3��-�O���������S=���,Ď�?Ӎu�8�ݝ�-�8���ɠ}��.��5Y� ��S�TR�T��Ą&'S�6����i�;�^__J�e���!`�rɯ�:���1         ���o��r�,�3v q��};Kz��E���o�:#�Hv�K;ǽ^|vY�M�+�A_[���R[!����y7Xw9�޵�X��Ο	�p6׹ӹFڤ �����驖����z��olLu��St`K1������N         DS�L?5�y��)�*v ��t涂�uZI��*&tf �3]�^p���,����kA_��t�B�|˔��t7V�^�]���^J��3]8��������`08�T.�U.�5�f�[�dWC����(���c��[�F'�Dr<A        ��V�������tq�8 zgz4��w��E͔)�<��Y{�����4/�����m}��V�e����ug�{w��+��]MIŮ�7 F����ؤ���� N\��j6�j4��β�k�����(��
l*&����js�o��         �]�o:?S��N�;��)&^�v���%�=C��pʂ��U�]G2}c��v��&ؚ�j����NW&����ޝR{���#�i߶�g3�3�+��`H%I���q���kj2չ;�Z��t�b��T-�x�=�2��r;         �HG殿w�����B~й�3�تv���%=�D�� í�M�.�YP
��6�;��z��v{Lv�0Սe�Rp���k8���3�3�)�_8��8�� �J��J��&&��O����=���Z�{eLu��y��9?W���A         �AT;t�Ϸ���H��bgp�Ӆ��z��%�=C���T�҅;L�(*����h���>�*����"78w����(�s�r]�=׾m�J	�N ���^�����T�3gzA��{jNwULu�������+��         dչ�q���[cgpbvNt�ޒ��'���l!�3훕���|ZQ_Y�ݿ��VCTv6ݍe�Rp�޶����I�;�)�_�=�h�R;���P(hrrR�>�ҳ�4���\_�t߲����2�o��@���c'         ����9���������y�oGQ�sfIg1� T.H�����=%��Gt��\w���r*�;����2])���m��o�>��.ޞi�De ��S�\V�\��d��v6T]m��U���
jd�x$�U�~X�ʀ?S         �?�n���b��d�Ď�a�D�>���Q��Ȁ ���3�.;���fI��P�;ʴ��J8��9W��:])���3��M+J϶��������qt�����v�4��Ӛ��f���h��ѱ@l&-&ő��o}�J�,         �0Y�������q�}N�d�<�V�w����-��yz� p¦��K�I��s=�V��| ӗ�j���ю1��ܝ¬)�#M�s�r=}G�}�r%<��S���ؘ���45���=����'��R""0�%���[�}O�(         �0Z<t�?︪�#�'$%�� [�s�;F�³�:c�A� p�N�0���D߿oT�\��|�������Y�\f68wsn[��������_�#�hap���fP*�T*�41���ن��-}y���jAi;�u���v������         ����[g�Wnt
�*J��%{Jz�9EM��Z ��t�t�LQͧ�Յ���;�R��=G�~����:]9q쒫��szZ7�:A:�ǝ�o����8}Ҿ��A] �3�{�J%MO���i��[Kr���Z9/>��r��U�;         �4�����|�dϊ��̦ˉ^t��^�̲.�U�H�~	 �Z�K{&�^xV�ѿ9<��Ω�L�da�_�,m����^:���]����n��$ڒ:����Ço��L����>� ��S�\V�\��TK�����2�ӑ�(b7    IDAT�M^� �f���6�࿎�         �L&z�꨻X����l6{&�z�9%]�+M ��9����?U��sz�G�ݮ#k��Y�m
�岬+�џ`��t�]y�u݇�Y�3��֣9g_��>�B�?�/o;|��~�7�"I_�ž ��e�����]h럎��:/O�n0�[��?��+Gbg         6����3���퉝�Ι-��t��& '"H�����_��u9M����o�<=���?&���܍�6ʺ2�]Ҷ.�sԚ��l�;������}����9�� S�P��Ԕ�5�k߮��Gݷ�cG���{^wx�r;         ���ʷw��r�>#���y�a�Ӿ�E}�9#:m� of��t��W.|�J�Q��v\��/Us��Ph�ukc'�t�9��/~��Ic]���������.���O��s��ζ �S�$�&&&t������Ѓ�}�׽��B�p�p19����          �ّ�>����,�p�,�0���{��޳��6� D D�糶p��J�_m��#�I{��-K߮�}�����-\\��橬ѕ��I�S��-'�*飇o~�_���T*%I/;�} =����ؘ����-Yj�2}�Z��� 3�[���9v         `+X8t���^Uy��m�� ��{�Kv���J�.3� �	_��˒~[�oo�o?_y���?���>Ս�Q�<�?{T��z*�����b;�=|�;�;�r�$MMM�H��S� ��9��e��{F��hLo~F�g�̔��x��w�і���w���]-=XT�# }�"��51AA��c<)-�x�j��Z�C��kNr���p\8��hc�����{Q��F���f����D��ݬ�޹���>V��>����6�?���K�yC�      ��L�����\}�t��fU�	ƫ�6/8fH�`~X�q�ƣfr���x��'>�_^���jp�?Gc蛳��w�ι�ޅ�9E�g`�ޕ">q�ͯ�XDʳ��n��Mɍ��)�?ix8�Y�3N�{��Os|cK3ڳ��s��ݻw����.�      �/����j�pw#��"V��u1Ш�����kc�R;��SUչ�^�o[�������w_yjx:�w�c�7���[�Sn�+��_�<�����>�r{DDJ��r= �744�"~󨱸�v�w�Fw���i[s0^��co�(      �{?Һ/��#���@iͪ���?z�X<��!�v�y*�t�\�xd�{sh�Ս�%����]3\5缀}�w�}^����������v���} >њ��G��mo�kpp��BA�rv��[����N|��ftJ�2rj^��k��t      X��yΛ_�I�,�JH)ű�obc;��uɒ%{]~�廻vb�U������w����ψ���Fg�OW?�鿸k.c�ܐ���]��iG��%�������W�z��<;������8p���{ٮ8~����{r|{�sz��;�u��      P�߱��z^��ȝ?*���J)�� �>t(�)�,$K|��3#�S];���������^����ij�k�ԮK��{����f5����;c�`��"����6����7�jr��>�n���>c�~����q���?	Ew����<#�16�N      <b������zr��9��@o�8b��8簁�k̾Y����:��+�������FīW^t�Սm;.�w�6ڻ����9���|�T4n�����}�Vg��M�o�i }444�����Ll��q?��(�T}'�zI���׿�      ��h�:��j]��_H�Jǁ^8t��8����w��v��,��[���3&�v��#���j�g�-{~~x���z漻;]��GG�7K� ��v��߿������nWtg�i[c0=����Z:
      �g{�N�Լ;>�)��e�%�8爡8dE�t ��]UվW\q�d� 31ۂ� @��OZ�0����K'�nH�\U�)�     @�m�p�Q�WGD.��j�h3~���x���� �K���<�t��Rp��RJ1::��<.>�O?���S��j���/      xb�o���ݥs�l�6⷏�?8s4��G�`��w��yUp�{�;�,���K)Œ�8��eq�U��;��]"rT�8=_[:      0}g�k#�(�f�Q�8u�p\���8��fT�t" 
���fj^ݶ�����"�S�s P^�ݎ{x(��G��֤'���釻w�:u���>Q:      03�?�m�슝_J��T:<�#��s��eå� P�F�u��}�t��o�o�U:  ��h4��������c��\:<��᪙�Sn     ��駛�xJ�EN;Jg��r�����x���� <Z�ݞW��Vp?�t  �e`` �<pY\x�p<��v,Pt�~RJ����R�      ��MlZ�O��ה��j�p�۱�q�)#q���V	�O�{��jGę�s POCCCq��q٩����10o�p,t95޻eӆ���      ��䦷�YD���s@DD�������g��S�o��@�=;�J���yS�FDxq
 �)��#q�Q���8|y�t$��+�זN      tϒ��U9������v�>C�O�s�fc��(g�o���!�k��SJ�� ��PUU��x��	K�G�X>�KGbQ���4����y���I      ����'Z;���H������=ֈO�?ˇ���v�����k��s��*�����l�q��ť���������1��4�S��[[w��      t߃�����^^-N_5S<��x�c�z� 3WUռ�bϋG�6nܸ��hLFD�t 槜s������N�][���y�ͫؼ���9      ��Z��7�%E�M�s���P<눡ў`n<����:���k��޼x����g�r; s�R�V�������|(��ĂU}@�      ����7�T�^:�^c����x�����ew�u�ɥCL�|)�ϛ�� �[�шc��4.;u8�vP'�ŝ�y#���KJ�       �%��qa��;���p6R<��x�cq�r� ��٥LǼ����誑�8��eq�	�8x�m�tC��48���?��V:	      �?��[?�"Ώ�.���������*�N�B�R:�t���-�mo{�^�����<)�0�LMM���=>��"�]:�T����ۆ��t      ��}���WvR�/K�`~Z:\�o5���(�,��}```�ڵkw���xj_xṽ� �_�f3N\�4^q�P��o��OQCջ��     `q���Q�u��?�0�:cL����9�NMM�Y:����g� ��0>:�9vi�wl#��N����41W�N      �71��T:����f\t�x����jZ�@t:��w�k_pO)�S: �GUUq��c���G��6wW����L���v��      ��-�]�j��9��Q���R��j8^y�H���> ���ͮuo��ۿ�������s�M|kW��p�o��:)�nټ���I      �zY��7��r�戬�̣�5ֈ�3-�� �쬪j�W\�p� ���w�F���3 �x����F����'�z�4�՟*�      {2�i��s��J�>U���W�1��@iC�v���!O�NG����qΑ�q�Ƀ��X.�Z�>6�y���)      ���<#�̩�T�����f\v�x<�����@������Z�SJ���`�H)�+���S��7V����^ʑ�i���i      ౵Z��=𒈸�t�hT)�:t$.;}4��l�>rε�h���y�M7�k׮{��X��}pG�ݿ�os�ZLr�]Q�3y���-�      ��~�[��c꣑r�t�g���x��C�lD� �Zڱm۶�VkG� {R����w�>;������ǅ���9�T��/&��F�      ��-w��9�?)���jV�ܣG����������SK�x,����}�= 4��8������8`�tz����7�N      �?�w�K�js���A˚�3��ăJG�'�R�mW������_ ��}��E���%�Y��更헔N      �W)�޵��qW�$t_U�8�������X>�9 ��P�e䵼��p�+;���Q�> ���'w�m��#�Y�[,��cg������JG      淽^��b�ԧ"�P�,tǊ�F��ؑ8h�� �KJi�֭[W�Z�]����Z�U���3��� ��<i�P����8q�#5�)�      �0q���w��s��0�<}L��y)�<�dɒ�K�ؓZ�YSJ�]y Odh��9f<~���(��9�Շ&6oxO�      �����6�H�J�`�F�������@�t ��N�S��v-�qv�  0)�8j��x��q�J��磜�t��/-�      Xxv��uI��Q����{��9G���������v��w��˚��DD�  B�9�|�����MŮv�4LK��1�|�ĭ�?_:
      �0�|��<-:��L�Kg�6�8���8m�W���lݶm��V�5U:�/���F�qV(������U�q���q�x�-cOR\��      �����~6��U:Ol�%�x��c�� ,DK���O*�Wծ�^U�3Jg �^�{�`����8kU��+T�%Շ'6���K�       ��Mޞ��\:{V�g���N�����`�:�t�_U��{���3 @�4�xƑK�%�Ÿ���N���qq�      ��{�΋s��K��і7⢓G����m`�cw�V��n�i("N-� z�}����ơ+�\9v�Ըprs�祣       ��֏�}��r�ݥ�������>OZ�( z.�d���ٱcǩ1\: ���P3^|�x���j���T]3�i�?��      ,>�m^����ͥs,v)�8��xɉ#1:��| �����#J��e�*���	  襪J���F�'����˩n���zW�      ��5���o�)�Q:�b56XŅ'��3���{ ��u��Vpz� P�ꕃ���b��Zݚ����t      `�Kyw#]�#�]:�bs�ʁxՙcq�
���8UUU�wm��9�O-� J�ₓ���C�s�^�r�j�t��>��Y�(       [ommiF��i�t�� �g����4�ֶ�x�k���Q:�#�,YrLD\U: ��R��Wē�������.�h�K՛�ln�M�       �x�w�h��sS�KgY���F����� �׹����~���Q��Q��? ��f��x��c�zy�n�L��ؼ��c       ����cC����9�5+�Ug�������"��C<�6w�sm�R �Ƈ��ऱ8{M�>7�"G����)��      �kZ�Nj\Q�_:�B�R�3W�'��蠽� ��RJ��rצ/W�� ���J���F��c�Y:�B�:UU]6q۵?.�      �L�v�#w.����`l��4�>�� �Gg���Zܫ�������I� Pg?����O�uJG��rT���ZW:      �t����{"w�S��فK�q���1>T�}� PG��m۶��jm/�w쪪j����Z:҈��:'�(e��9�29W��      0]c��՗K瘯�;`0.:eD� ����%K�("�&����Kg ���٨�9ǌ�o9�Z��e>�~�h�8ni�*�      `�ni�F.�����2�TU�s��3��� 0M�XZ^��{��i�3 �|r��x��#16���"��ۛ�S:      �Lm����JU���9�с*.<i4N}R�t �WrεXZ^�w�7�t:��E�`�, 0�<�������w[�t�zK��Llj]\:      �\����-�鼨t�:�I3�;~$����|��m۶��j��Ҋop�t:��r; �ʲ�*.9u,��o�t��J�w�����1       �*w�9��K稫��KNUn��[�lٲ�J�(^p�9?�t �Ϛ��{�H<���f��;�Q]t�'Z�JG      ���ͭ�Gn�,��]:K����G����F�F �o�N�x����<�tf� ���z(�?q$��j�ȍ�ډ[��t      �n��c��"5�Z:G]�T�ғ��7KG���ˋ�#�� `�8t��x��c��xn������7���1       �mr��?�\�Y:Gi{�5�姍���#�.*�������_��  ��*.9e4�ާQ:J19b"�͋#R.�      ��R�f��iK�$���@\v�h,�s �c��w,+�h�=�T�� �@��>e4�Z3��G���z��m���t      �^����W�Z[:G���♇��yǏ�@c~# �W5��Ӌ(9<��Ԓ�`!K)�3�7�����>W�_Nln}�t      �^۲i��"US:G�4�x�q#����� �BW��]����� ���`\x�h�.��{��3\��J�       �j{�:"�W:G��T�ғG��}��� �bpf��Śn7�t�Ю]����R `1ypG'n��ñ�v�(=�#�J��Y���|�,       ���3#w>�R,���+G�Gb�H�}� �h�l۶m{�Z�N������w�>%���o�Wqɩ��f����R�Rn      ��ͭ�T��t�^8xE3.=mT� �k���������真Zj6 ,VC�/9q$N8p�t���Q}rb��w��      P�����gJ����N��f* ��]��Yp6 ,ZU�xޓ�㙇���9�h7_�r�,       ŴZ�Nj^�#��t��Jq�!��c��Q)�@	)�b]ow X���f0~���h��5R�?M~����      P��6]����xM�sѬ����F��.�7��<T��]��o��v�}O�� ����`;��W��C����\�?w�^^:      @�����ˑ/(�c�F����Gcղy�� ������׼�5��=�ȿ���%� ���e��䔱X12��AN߭v���      P7�H��H?,�c&V�6��S���F=��I%����i�� {�|���N��+���LW������Vߟ      ���ͭ�Gn\9M��2�V4����b�|[� \UU��[bhD�� �mx����8��7P:�4T�ۼ�3�S       ����?��]�s<�����8��f ,*E������sNqJ�� O�Q����F�����8җ&ƏY_:      @�M���7樾\:�c9u�P����hT�t `ϊ,5o�{�ҥK�����= ���+�1�H��ɺ���z87;�{�|o�$       ���/v��|�gS��"r�^�}�������| ���{�{>�я>�ϡ}����� �̜�z0~���EN�i��7N���o��      0_<�i��:�j���c��<�~�!���  ӐR:��3K�O+0 ���n�Yj�FD_��۳�&7o���)       �6�靑�;K爨N�:�)4>Z:	 0=)��/7�{�=�� �C��n���o������
�#�/�H�T      ��+��@\�s<X*A��`���'6�>XU��J�  f�D��������qb?g ��񫯾�����6������o�~R"HjT���ܺ��l      ����[[wU��k��龪�����wFDLMM} ".� ����������>%"F�9 ���ң����C�|-7�̈�[��Q�<q[����L      ��h�m�6��@_���ݩ��[n������zk�yS_s  ��R���o\�ϙ}-�7���� feWJ郿���ںk�9~VD��=]�}�Ow�Q��s�    IDATf      ,|�;��~�ʩ����Y������UU��=] �O���k����Pp�y ����+������s��T��̈�=NѩR��[?�Ɖ��      X<~�w�ɪ��srT�ɻ�~��������n�z{D<�� @w�n�=�|z?� ���O��KkۊX���Շz� ����Mo��g�      ,R[n��)���݄��������,��Z��ko ����[��hD<�_� �Y{�����D���;'Όߏ����G��32����?      ����FzmD|��禔�r�xQ���5��?��5 �RJ��Z�����6hll섈h�k 0;)�]u�UM�íVgbs�9һ���su�ݷ\�p�      ���skk{�/��v���Uu��Mo��h�:����m�>�vk> �3�###G�kX�
�qJg �7�'�'7�y]��-��Su���?׍�       xl��q�sTޝӪ��������Vk*"�ߝ� @/5���5�o��R��P ��=�u�֏����ͭ9��8��+��7��       �ie��&r�׹���Ӊͭkfy񌗰 E�m�y?7�+�@ͥ��{���5��'7oxk��ED��9��4P]���kw�v>       3���kw�@㒜c�,.ϑo�ؼ���ο��+??��� @�,��Vk8"���, `N��d��ۯ}WU�6"ufr]J��|�����      `f&n]����fxY����6�}.�SJ9"n�� @_��sN�ԗ�����S"b�� �Y�oժU���A����?���ў���'��[�1      �����7圾:͏��j��6mxg7fWUuK7� zjٍ7�xX?�����i 0K)�����,�?��7����j��%�iWjƥqKkW�f      0C_�����tq����l��x������n�^�n�SJwu�< �7������ӗ�{J�/ `�r������~�_WU�9���ӟn����n�      `f��p�9U�9MEռl���͹)��s�P7� �/�ԗ��6� [�m�vg/����D�.��S��K����i/�      0s�gě#W��W=�؝�ꒉ���M/榔��� 躅����j朏�� `Nno�Z;zu����3R�pnv.�[�o�j.       3�juR5xqD���/�H���E[6mx_�ƮZ����W� ]qJ�9�zH���E�P��  ��s�����6|(�ꅏ�O�NTo�������\       ff˦7~;R�'�����λ����r���ߎ��z9 ���_��^�y�=�tJ�g  s�shh�~��c��E�~'ru��w���L       fn���1��X��y[6��R<O)�|9 07UU����^H)�� ��߯]����6qǆ�E��)�k&       3�ju&"�ѿ�v�n��������_3�;%"���=��'�a 0K9���r;      @�����V��#���~� f������ӂ��7��H)=��3 �9��o-       ""RJ(� xl)�{=�����눜�h/g  ��R��������       SSS�EĮ�9 �Ǵ������z9����s�� ���=�      @m\s�5��>Q: �ئ��z��i�=�tB/� ��h|�t       �e��@���#�ӂ{�8< 0'_^�n��K�       �_�l6?��9 �=��tw X�<�      @��u��7"��t `�r�'�����o��}"��^� �MUU
�       �R��w� P_G�Z��^޳��Ν;mo����W\��!       `O���; �Wc||��^޳�{JI� jʓ�       ��W\�݈�F� �c�YW�g���: ����6��        �'缹t `�z��w X|�t�       ����z��'�V�5G��l `�>�v�ڝ�C       ��y衇>[K�  ����s���=)�/Y��؈��� ��y�      ��k�Z�RJ/� أ��|�;���=)�眏�Ź ��5�;Jg       ���9o*� س��N�ɹ�8T� j�_֭[���!       `:��; ��q�8�'���z ��ͥ       �t]}��wG�7J�  �h��s�O�Ź �ܤ��      �Wrξ��z�Ig���n�aeD��s�9{h``�ӥC       �)�@=q�7�t��^lp�� ��ck׮�Y:       ��ҥK?�� ������Q�>���v��� ��v       ��/�|wD�Y: �몪�zw�܏��� �5����        �d� �S׻�]/�WU�� 5�s��u�_:       �F����t ��r��.��S���n�	 t�'�      ������#��s  ��RzJ���j�}�ƍ�"by7� �B�      ���w� P?�n��Ʈ�ǻZp���y `��T�       0)%w ��v���yW�9gw ����]�vg�       0��㟎���s  ��RzJ7��v���� ���9�}�       0W�_~���d� ��圏��y]-���lp��i4w��        ݐR�x� ������o��Gu�< �+�[�n��K�       �.�� ꧞����C"b�[� ]qgJ)�       ݰu�֯DĖ�9 �G���|��:�k���1�: 莔�'�      X0Z�V'">Y: �h�F���:�k�N�ӵP @�(�      ���} 5��e�]+�����^���+�]:       tSJ��3  ��s�����Z� 芏�        �v�W~3"~Z: �(����sNqt7� ��+�       X�RJ9"|' �R���ƍWEĒn� tG����<       ��o P;���o_э��Rpo6�O��9 @�|oݺu?,       z!���� �G�J��+���Jy �+<�      ����7��{���9 ���s�J��+���� P#^�      �"��� ���s�� سN���       ��RJ��@��g�{���n� �]���W_}�=�s       @/MMM�}� �����w��]�E�^]� tAJ��3       @����o�� �B�y�ƍ����9�;���� P#^�      �"b	 �Gj4G���n܏�� @���?�       }��� �G����9�s�
� P�z��_��t       臩��ϔ�  <J��)%w ��ϖ        �r�5��?*� �ws�Ϲ�ލ @w��      Xl|W �Q���j�#b�\C  ݑR��5       ߕ@}�sNs9`N�e˖͹� t�ĕW^���!       ��:���; ���u�]w�\�S���n�y�< �5�M)��!       ��֬Y��Z: ��fsN�9�s�
� P�-        �����oG��,� ���v��TpO))�@}(�      �(�}g 51׎�\�G��z �kvo۶��C       @	)�ϔ�  �B��s t͗Z����!       ������ED�t  ""��o�ᆕ��\� ݑs�$:       ��ڵk�(� ����o�ᆑ�^<�{�ݶ� j���ϖ�        %Y �QE��s�xVRJG��Z �����>W:       �d9 �G�y�]�Y�c�z ��~p��W�S:       ���tlp���t:���
� P^�       W]u�"�ǥs  UU6�k�0w�C���5       �w�+  ��9�� �U����9       ��%q PG���Y������+f; 莔���۷�t       ��ϗ  DD�A7�p��l.�U�}``��v ��n�ZS�C       @l۶�K�{t (/����fs�
�)%w ����Jg       ��h�Z�#⛥s  ��Ϫ��j� ݕRRp      �G�]: �@_�9gw ��      ��RJ_,� ��t:�+�϶M t��m۶}�t       ��N�cY �@_7�G��; ���V��)       �䡇�JD�.� �]�|���n�iiD�;�a @��=q       ���j툈��� ĪV�5<Ӌf\p߱c��� P_,        �(�di �W-[��_4���Й^ t_�Y�       ��[��:��a3�f����[� @�=x�UW}�t       �)K� �:�Κ�^3�{Ji�L� ���)�\:       �ђ%K�;J�  b����#b�,� �˫�       �1\~��#�k�s �b�RZ3�k�`~�*5       x|�/  ���^3������ �F�a�;       <����q PX�7��t�M�DĒ� �j˺u�~X:       �Y�ӱ< ��{�ƍ3�Ϩ�k׮53� t]���       �V�^���x�t X쪪Z=����� t_J�K�3       @ݝ����Z� ��UU�fF��ɇs·�( �u9篔�        �����N��f&��Q�=�d�; �R�j�       0TUe�; �7���
��f�� �kǶm۾[:       ��v�9 (,��f&�Wp����Vk�t       �:��W#"�� �Y�y�L>?ӂ��3�< �]^�       �t�5�<w�� �Y�6�_��{GĒ� �(���       3��� `��{�ƍ��O��^U՚Y� ���^�       LS��w� PXUU�����~��鬙U ����       3PU���@a3Y�>�{Jiڇ =q�UW]u_�       0�TUe� 6�e��.�GĴ�� =�n       ���:���p� ��M��>�{�yͬ�  ݢ�       3t���#�_J� ��,��f�����i
 ���J  ���Ǯ�>���6g�CR%[�\�
I�6E��.�m��A����.�`A�ݹ�@S&��WзiP�v
[�*�rdQ_4CΜ�za����e�:�����9$�;ba=��     ��r� ������< <z�8:l      ��Lw� ��#_p��7�O<` ��m��g^�       `�� &O�>P�@�R��* ��y6�m�       �hmm���  S������|�@�q� �ƫ�       ��:u꣈��w ���|���|�@��<�? ��Tp      ������; L�A;�*�GĿ~�$ �C����        ���; �Uk��A�w���A�1 �p�����       `�e�O{g ��;���Aܟ�  ���:y���{�       �%g\ :��u�Zp��Cd ��^z饭�!       `��Z�����}�gϞ]��g: ��      �!���+��� ��w�yg��K�ܷ����h�  H�       ���  6���_��K��K)�� Gf:\      ��ad :�a�n���Z�w ���       #s ����3ӂ; tt��u�k       x2�� tt�n�w Xl�����       �	w �� �t� ���      ��|���#�Z� 0a��~� 84
�       ���f���Y� 0a����< p8j�?�       3�� ��Z���k�
� ��0�       �h���N2s�n���7�x㙈8�� �e>�[p      �G(3��@?O�;w��^_سྲ���< ph6�^��^�       �8����� `�677�\q߳�>þ� �����l6�       ���|�����s ���9¾g�}>�[p�~~�;        <n^}�����9 `�����_y�Y ���z       �ǔ;y �d�/��Z��h�  ��?�       S?�  �����=��/3sϿ �Z��4       �s ��C-�g� 8<��\�       ��9 �g�����Z��; �������!       �q�����+��f�#��#� ����l6{�       ��Q)E� ���l6۵Ǿ�/�x≯��{ ��d�W�      �!y��/D���9 `���<yr�!��
�{N� �ǫ�       �p��~�_��kW]� �8����        ��Z��9 �$3��^k���� �!       ��y ��
�{�% �p��5h       p�j��������w-�����É �^�t���!       �1g� :y�ww ����l�Y�       �8�Lw ��wv�Ů��x��  �s�      �C�����{� ��z����	 8<�֟��        ��_|q��� �����ZkF�- ��R��;       4Pk��u �����z뭧"b���  ���       md��; �q|6���;��qܵ .�g       h#3��@'O=�Ԏ�������Í �f{{��3       ����n� 0U�u�w,�g�w �����Ƈ�C       ���{g ����|����� }|0����!       `
�����3 ����^k�q� 8\�VO�      @#?��>����9 `�2s�����ݾ ���d8       4��5">� �h�Q���w�{ �w       h�]= ��cg}ǂ{DXp�>�      �-o[�>��n� :��*�      @C������q�]� �0�
      ������-��Z3"�p�q �{d�C3       4���� �����x�g"�ȡ� �v�������!       `b��@ko����w�������Mx ��y"       [__w_ �lnn>{���)����{� �Z�'�      ���~��W"��9 `�2�q�{
�a� :�LO�      @F� �w X`�       ЇQ: � 3���g��w� Є�;       tPkug }��^kUp�2���       Ї�; tp��ء ��tX      ���@7�/�G� ����       `�J)��  STk=Ђ��d �t��_��       �h{{�W�3 �D��S 8t�        SUkuo }�]p��ff>�. p��2       t�ꫯ^��+�s �}���Qp?}���14� DDD�ի�       �/�t ���ٳg�?��;
�kkkO�� DDd���       ���= ����uG����˓m�  ��)p       �֪� ����^p���; t��       ݹ���qܽ�^kUp��      �/w� �Gf�����/�6�qtH      ��J)�����G�-����~�;       L�w �cς{DXp��6^{�O{�       �)Sp�>J){�-�@{�       ���֖�{ �㎑v� �Yf:       @g��������; LM�u���	 >�8      ��2�f�{� �	ڽ���
� О�;       , #u �����{��d  �}�;        F� �� �H<�       ��> t�{�="�j ��̴�       ���� ����[��gϮG�z�8 0q�8��w        ���Q� 0A'f�����
�yr�� �i����        Dd��; t��3�<u�Ϸ
�����>q `�677�      `d�;| �`kk�V��V�}Gw h��l6��w        bG� ����H5R:    IDAT
�y�O �4O~      ��X]]Up��a���^J�� ��Z�      `A|��_�c� 05;.���h� �Lw       X/���<">� �&3ou�-�@_��        ���: h��j� A�ա       ���@{;�3ӂ; �g�       ��| h,3o�����\� �s(      ��m� �ގ��D�, 0i^k       �E� ���7������� .�       �X��@c
� � �󹧾      `�x; �WkUp�E����P       �ł; ��� `~�ҥ��C        ���h� �Sp���l6{�        n�A� ڻ��~�����X� �Ɂ       ��˗��@{�f�Y��Qp��ώ�� ��q�        ��f��fD\� &&��׏G�(����D�< 0Iz        vt�w  �����7
}� �$9      �b��w  ��������|�� �9      ��Lw� �����Tp��,�      ���*�@c�����8*�@{�       ����@cw�-�@{^g       �ɝ> �ws����|�c ����        ���*�@c7G�KDD�Ղ; 46���      `1�����Xp��v �)�8      ��Lw� ���q�c ���|~�w       �^�8*�@{�#,�@7+++�       ���� ڻc��֪� m]{��7z�        �� ��촗���-a       XP[[[���=� ����       ��=zT� ڻ]p�Lw h�A       ԩS��E�F� 01��7?  m�Z�      `�y;; �u<B� �(�8      �b3^ �Z-�@/�      `�e��} h(3�(�� &'3/��        ����� �����A `rj�
�       ��.�  S��ke6���8�9 L��;       ,��Tp��j��-�G���Y `��      `����n �f�ّ�����;	 L�C0       ,6w� �������0
� �X��R�       ��J)������������ �e���      `����n �a���󣽃 �9      ��� ��Zp���C0       ,6�u ��Z�Lw h�!       �|>w� �mmm���Pp��������!       ������ ��0GK��h�  01Wf���;       ��R�w h,3-�@�       ����w hlǣ%3��-`       Xp���� ���\+�֣�� ��8       ��;u�Ե���; L�Z�� Ж�;       ,w� �P��h�Lw h�R�        ������,�@��      ���� �̵Rk=�; L��/       ,��t� �Z��R�j�  01Wz        �Wku� mYp��2��       ���;  L�Z����) `J�qTp      �%Pku� m-��� e���      `	xK; 4�Vj�G{� �)q�      ��a� �Z+a� �Q�       �@��? �uT� +�8�      ��v hn�d��; 4d�       ���� `b�J��H� 01�       �j�F� ���J�u� �d�_       X�� ��%3�����m�_       X����D��; 4�����       K��z�w ���J�U� �v횂;       ,�R�;~ h��:��Tp���~�i�_       X�8�����
� ����^zi�w       `�֫�3 ��d�P"�� ��n       XG�q� �Z�Rk�� �8�      ���L� ��P2S� �Qp      �%q��%�� �V)�� �x�       ��l6ی�y� 0�9��(�� ��l�        �w� �H��H��#�� ��l�        ܗk� ���C� 0!�       �\��@#��A� �L�^       X.�� ���JD��A `*j�
�       �\��@;���Z���      `�x[; 4�� -9�      �r1f M)�@c�       �\��@;
� ИC/       ,� Д�; 4��       K$3��@;
� И�;       ,w hG� Z�T7       ,cv �NQp���qTp      �%Rku� �%"J� 0!��      �%�m� Д�; �TJQp      ��� ���w
 ��q=�       ��]? �S���R�C/       ,� �Hf�c�  0�V�^       X.����Z�h� ��       �%3��@;��%�       �\�qTp�v�w hK�       �Hf^� &d�� ���;       pp�Vw� Ўw hI�       �K)�]? �c� ZZ]]u�      �%2���� `B,�@Kׯ_w�      �%2�1; h��Z-�@Ckkk�       �Dj������K�Ղ; 42��C/       ,��|�m� �N-��� �lmm)�      ���]? �SKD��S �T���{�       ��w hj,a� �pႧ�      `�9r�]? �c� g���w      `���� �T� Ў/       ,�a���  2�̴$ m8�      ���� M�Rk�� m8�      ���� M���w       X2����D�w hÁ       ���֖�~ hǂ; 4�e       �d�����@;Ղ; ��n       X2.\p� ���^       X2��l��y� 0��Z��w       XN�{ ��Kfz� ���        x �d����d��      �rr� ml+�@#ޚ       K�[������
� �@�U�       ��; hf��Z��Os      ���v hf�D��; �1�        <�v ��v	��@+Gz        �j�  0�V� ��z�        �q� �R�J�U� �p�      ��t�w  ��q�Kf*�@
�       �d�y�!"Vz� �)�̭
� І�;       ,���{�z; 4Rk�.q�w �^       X2�i� )�l���� � 3���        �w h�ֺ�� ��Z��f3+�       �D���zg �	�(��; LœO>��       Kdw� Ўw h�S�       �\�qt� ��Z���R�C/       ,w� �Nfn���� �����       K�]? �������t�      �%� ��Pp����;        pp���q-�@K�8>�;       p_��;  LEfn�q7{�����;       p_���R�f����� ��(�      ����f(�@3�8^)�0\� &���       �������X� �b�+e>�+�@;O�;w�D�       ��2ӛ���#G�\)�y�w �����.      ��� moo_)W�\�� ���|�       ��<�;  L���ǯ��l�[�� �T��B�       ���q��� `BƏ>��r��ծQ `Bj���;       ����F� 0!Wg��x��~�k ��_       X�;  Lȕ��Qk��7 L��;       ,��lv$"^� &�v�=3-�@;�{�����!       ��;v셈X� &�v��� ���+W�x�       �0��; L�Ո��K� �}�w        `w��?� &�b���ŎA `r�      `����>��]p��c ��?�        �]f�I� 0%��I�w �"3�]�       ��j�YkUp��j�#n�o~  ڨ������Wz�        ���[o�O�� S���F�(�ߜs �Y�z��7z�        ���� ��8�������|�0       ���o{g ��)�\�Pp�n2S�       �;} h�f��DDd�'}� �$9      ���Zp��J)�F�(���h� �s      �s�ܹ�B� 05[[[��� ��WΞ=�\�       �m׮]���ѭ �Y[[�q�?�W^y�jD\� &hǿ�       �m>���� `�������;�2��S �2w       X �w� �ާ/���Vĝ��t
 �Uku(      �Rk��� `�n��+�@G����lv�w        ����_���z� �	��eWp���?~��z�        "�a�� }�[p��*�@�;        ���� �(J)�       � j�����Z��7�|������u �0�Z��;       L����W2�s �}��n� ���3g��N�       0e�.]�fD� &�V�]� ��Rʷ{�       ����� `��`��Z��w       ���tw �(���qH      �N�y�!"�c� 0U�0|t�Ϸ
�FD� �����_�       ������ӈx�w �����o��V��ԩS�"��.� �\YY�O�C       �e�7�@?�^{�7?��~�a  ]8,      @7�;  Lؿdf��A� ��;       �7��J��۽s �T�Z���
� � j����o?�;       Lɉ'�,"�� �*3���]p�u  ��k׮���!       `J2�ozg �)�����w ��̿�       ��֪� ����� ����       �T�>}����V� 0e{.�g��; ��ܛo��G�C       ��R�KD��� SVkUp�E��g       �Ff�������Qp/�(�@g�       Ќ;z �lς���~���j� �Cf���o���;       <�Μ9�BD�^� 0u�8����(��f�1"��@G��c׮]�v�       �8+���� ����+�\���_��Q `����       g�����  ��]ߩ���~ 4Tk��3       ���ܹs'"�?�� ��]����������9s���       ����������s  (���% ������       �1��� ��Z����� t�0       ��l6+�w�s  �����8~�& ��?�я~���!       �qr�رoEėz�  ""b����ʊw X%3��w       x����� � ���=���܇a�eD�&� �=�R�      ���zg  ~��ѣ�/��:u�Z��7m" ���gϮ�       ���g��^f�a� @DD\����wOo���{DDf��y ���Z����w�s       ��`�� ���̬w�pǂ{��� 8(�k       x2���  ���N?ܱ�ۗ�.�s�����!       `��9s�Z�� ���Tp�%ubǿ�       �܋��C  ���^J�šF ��?�        ���;��������ꢛtUEIL�"(��yf�g��a�e�	K�^�0��#������cB@6�� �YT`�e�Q��FԤ;KwW���c��z��s�����oչ�O���|�I�RzZ� �[x� &���V:       &Q�۽OD<�t �ORJ���8q�#� �j~~~�q�#       `�|�=��  �ɚ�]v�Mq�H� �5�9?�t       L����J7  �b�s���pʁ�I_M �N����m�#       `�,..^�RzH� �[|e�Ν'N����SJ_Y ��n߾��#       `����<#"R� �[�p�/����~ (#����       0a�Y:  �V9�/��k��眿0� `#�����]JG       �$�t:??Z� ��?�N;pO)��C @1ۖ���R:       &AJ��� �Bgڪ�v�^U��; ����       gW�u�RzF� �;�/��k���t�M�� ��z��KG       @������8�t pJk�����#�+#� 6��9���       �f9g! Z(�t�}��z���v��s>�2 (�9�       ����O.� |����SJ�t_?��=�d� ��n����       �F۷obD|W� ��θQ?���l �zv�        h��ҳJ7  ��s��~Ɓ��> ��Rz��C�fKw       @�t:�{F�ϔ�  N-������a ��{�|��O(       mRU�s#q �^���8q⯇� SJ���       �-r�)"�W� 8��`pƍ��_~�?D�ׇZ ��8p��JG       @�z�GF�E�; ��:~뭷�p�o8�����wH1 ��m���٥#       �r��: ��_�u�|�oX���sC� F ����b       6����s��zj� ������Y�9gw h��v�?]:       J:q�Ŀ�9�S� 8���Y��g��� �����W�       J�9?�t pV�}ff�� ��鋋�w)       %t�����(� �Y�y���n����<�" `T�<�^:       JH)�B� ��2p���xD�0�" `dr�/(�        �v�����xN� ��q߾}_;�7�u��s���{ �{`��yD�       ��o����]�; ��Z�&}U����; L���..�        c�� ��[��� 0]�������#       `:��#r�.� ��gW�M�����|fc- ��l=~���KG       �8�K� 0QV�I_��}yy�� &DJ��Çϔ�       �Qj��n�� ��䜇7p��+�_�P 09���~�t       ����m�# �U���/��j�qU��>�� `�RJ�       S���*"~�t �j�ݱc��j�q���Ҫ�� Z�g���}JG       �(���?!"�{q �k٢�z��s��; L��+�       L��`��� ���^U��Z_ P��<xp�t       Ӂ~(���� ��������`�����o���#       `�fffvGD*� �^UU�ޢ�z�w�ޯG���U �s�ź�W���       �f�~��#♥; �59v�ȑ/����:x[��� @+\4??���       0���?E��� ��|�����~��)�O�� ()�|I�       بC��F�ť; �5��Z�yM��� Z�ѽ^�A�#       `#�9�8�t �6kݠ����\[ �9��       �A/.  ��Z7�k��OF�`ME @<���ܳt       �G�4����(� �]UU���۷���� �6�:33��t       �Ӯ� �����ݻ����i��s^ӂ h����u]o+�       k������t �.kޞ�y��R2p��t����疎       ���"b�t �.���y��X� �����-�#       `5���{D�sJw  �s��Z?����̌�; L����J�       X����]��t �>)�5o��<p��K�&"n^�� �v�9_�sN�;       �L�����9�,� �� ����~h���RN)���x �5���W:       ��رcGo&��    IDAT�]Jw  ���}��ݲ��y�1��T< �*�K       ��,--mM)�b� `C>���k��X�� �v��n�a�#       �TN�8�܈�W� `�r��ڜ�k��RZך h�����       ��><�s�S� ؘ�n��5p?z��'#��z> �Ɠ�����       pG7�p�S"�� ��������Għ��Y �5����       �F�9UUui� `þ�w�ޯ����G���x �U���v�S:       ""�����\� ذ�������:�� Ze6"��;       ��s�/� ��X��|���`�w �)��5MsA�       6�^������� �ƥ�ֽ5_����[n���X^���֘��}�#       ���(  �����i#7M�x�F�  Z������.�����t       �O�4���w��  ��{���z?���OZ�� h��[�l�;       ��R�  `h6�1����c�< �9�_X\\�W�       6��i/� �G7���SJ� h�m+++^q      `�RJ��t 0<ݘoh�~�ȑ�Gĉ�� ���^q      `\z�ޣsΏ,� ���L��{]׷Għ6r �*�VVVv��       `s�9�R� `xRJ7^r�%_���GD�?��3 �VyQ�߿w�       �[��y\D<�t 0<�ؖox�zB h�;�KKG       0ݪ���� ������ 8���n�>�#       �N�n��D�CKw  �Պ�/���OG�э� �ʝRJ��t       ӧ��*��˥; ��lݺ��=d��;v���>��s ��������/      �t���{fD<�t 0t�]XX�y��lx�1����֙YYY�KG       0=:4^o��4�M�P�)��� �u����~�t       ��ȑ#Ϗ����  �/���㜡ܫ���a� �N�9�j�       &_]��"�%�; ����a2����]��_�Y @��\�4�*      �d���QD�W� �[�9��a4���I^q�)�Rzi�       &����r��Jw  #󑺮��q�0�CyR h���#;���Jw       0�n��}q�� �h���lXgm��R��� ڧ��n]����8       6����{EĞ� �H�����fgg?ǆu �:���{v�       &�������; ��ɳ��>�Æ6p_XX8��y @+�Z]�甎       `2,..�?"�[� ��ZXX��a6��{DD�yhO� �tﹹ���       L����&"���  F���<l����P� �V����޽t       ���v���Jw  �5��P�+++^p��7_U�KJG       �^9�RjJw  �7�;p���K��R�q�g �s����\T�      �v��z�."R� ��/���O����#"r�2�3�֙����JG       �>u]o��N 6����رce�g}��R�а� Z�i�^��#       h��������t 0zUU���������� 6��s�sN�;       h����e����  �#�����޽{?��� @+=���?�t       �u��:"�R� ��7�|�G�}���)�2�s����u}N�       �j��Gr�;Kw  �R�h]׷�ܡ�#"RJŹ @�䜿~~~W�       ��G�l� `<r�#ٌ�d�>�`s���/����       ���i��/� �O���Gq�H��{��#�Q� �O���-[���t       �W���"�S� ����̇Gq�H�;w�<>����zV�4?]:      �񚛛���  ��S�w���Q<��{DD��C�: h�W�u=��/       h�����qy� `�F�� ���l ��2??���       ������#��� �x��&o�~�-��YD�� @;�;KKK��      �)��t�)� �]����������[SJ�� @k����㗖�       `trΩ��_�n� ����%�\��Q>�.���Gy> �Z��t       �����]D�t� �����Q���G|> �Nۖ����       `����΍�N� ���>�>ҁ�֭[?��� ��RJ?����X�      ��:~��K#��Jw  E����`�����c�g�� h���v��KG       0�~��E�ť; �b�r�޽_�#���1� �P���#���       l\]��`08[J�  e��F���}0��&�R��4���       `c�o����xX� �����z���� ����Q:      �����ߝRzY� ����Ǐhԗ�|�^������ Z�1�nwG�       �'�܉����  �I)���_���g���F�= �n)����Kw       �6�~�'s���t PV����g,����� �ڽgff~�t       �w����`p(���* �^�3p?��>?�� �V��^����       ��7������ @q�WU���h,�;v��?0�� �Vےs�o9�T:      �3����N)�J� ��d��ݷ�㢱�٘���7�� �V��i�c�       �l0���8�t �
��Ec����3�� �vK)u����Kw       pj�^�)�� @;TU5}�ݻw�uD�͸� Z���U�#       �NKKK���t ��p�y�}b\��m��R�r h��6M��      Z����݈�W��oz�;V�u�X���� ���\\\�K�       ���i?_� h�����y�X�'N�x_D�y' �j�ZYYyi�       "�����+"R� �=��z�X��eW\q�7RJ�s�w �wq��yD�      ���رc/I)ݿt �*_صk��y�X�9�?�� @�UUU���N�C       6��i~8���t �:׍�����}' �z�����t      �fT�u�RzUDl-� �K�y���{�D�M� h���K��;      �1���{a���; �ֹ��[n���/��}�Ν'RJ��� @�m����'       �U�4Dį��  Z�u]�:�KKȮ/t/ �b9�Gn߾�E�;       6��sJ)�""�K�  �s��Ľ��E�a������N�sQ�      �i����S��q�; �v�9_W��"�={�|)">S�n ��r��TUuu]ץ~      `�-..^�s>P� h���߿��%..6�9���� @�=|���/*      0�r�i0����- @;圯-uwɁ���� گ��+;��E�;       �M�׻8���� @�]W��b�m۶�QD-u? �n9�s������b?�       L����#��; �V�e�֭*uy�����±���R� ��۷oQ�      �i�sN+++�����- @����ֻ��/�^[�~ �媪����\T�      `����D�cKw  �w]�ˋ�SJ\� h���9UU]]�u�_�      �X���术,� �����K�_t(�gϞ/E�'K6  ��۷oQ�      �I�sN+++�����- @���e�]vcɀ6����� @�UUue�����       ��i�G�cKw  �R��tC�{J�J7  �s>'���C�͖n      �����O)��t 0r�זn(>p?r�ȟE��Jw  �!7�|�KJG       L�C�ͮ���6"�\� �7����tD�{]׃��Kw  �!���^��S�;       ���ѣ�?Q� ��޹s����UU��t 01��_�����!       m��t�s�[� �(ו�h��}vv���8^� �����[:      ��<8WU��1S� ��-[���tDDK�7GćJw  �#��������       ms뭷�����  &��.�䒯���h��=""���� �dI)�rii�{Kw       �E�4OJ)=�t 0q~�t�7�f�e˖k""��  &�=�?���       mp����� X���~�t�7�f�k׮/F��,� L�'v��痎       ()眪�zeD|O� `����ݻ?]:�Z3p��H)�f� L��үw:��Jw       ��4�SJO(� L��������^� �H۫�zm]�[J�       �[��@UUJw  ����V=Rު��ɧ�?W� �H������       �T����`�Ɯ�9�[ ����]�v}�t��j��R��t 0�.�v��)      0.���K��� ��z{J)�������A��� &J�Rz}�ӹg�      �Qk��9�/� L��R�ۭ��ݻ�#�� �ĺGJ�59�T:      `Tz���q�t 0Ѿq�ȑ���v����rJ��; �ɕR��^�wI�      �Q��zK����ݥ[ �������KG|���#"�A랺 &΁n����       �6??�҈xx� `���Z��n����.����z� `�ͦ�ް��tn�      �a��z�<缷t 0�9r佥#N���;v�D�;Kw  �ǏE�      �a�v�w�9�!"fJ�  �꺾�tĩ�r��sn�� ��yz��{N�      ���9���oGĽJ�  �/��ڭvk�[�n�È8R� �|9��l��Kw       �W�����t 0����^W:�tZ;p_XX8�� �(�#�u]o+      �V�^�"�WKw  S�=7��8���#"rέ}� �8?>??�T:      `-����s�o��;�n �CJ���V��9�wE��; ��s��^����       �Q�uUU��DĽK�  Scevv���#Τ�����G#�}�; ��s��N��Jw       ��������Jw  S�CW:�LZ=p���9��	| `�l������ҹ�C       N���=:�tE� `�L�6�����;"b�t 0U.:~��+KG       �J��;?��战)� L����rM鈳i��}�޽_��?.� L�MӼ�t      ��u}���["�n�[ ����.����g����Io)  L�^��yD�      �o���k"⡥; ������1)��q�t 0uf��zS�4^>       ��v�;"�_� FaPU�[KG��D���������Jw  S���x��ÇgJ�       �W�ӹ(���� �����ݻ�\:b5&b�QU�D<� L���x㍗��       6�n������GĹ�[ ��s~s�՚������5q[� `j�M�<�t      ����^?Z� �Z'N�8����51�����#�Jw  Sk&"~���ܷt      �yt��}�� �T{�W\���51���T:  �jw�����nw{�      `��z�G��^V� �z������ѣG����Jw  S�)���S�      `z5MsA�����t 0�RJ����w~g鎵���{]׷G�5�; ����i���       �S�߿sJ��q��- �t�9��_�£�;�b��'M�� �dJ)��i��-�      L��s��9?�t 0�RJ������ѣG�_-� L�*"���t�[:      ��^o_D<�t �)�������#�j��u]/G�[Kw  ��]��z{���^:      �|�n�1�� ��Rz���±�k5q����`0qO� �)���S�      `r-..^�RzSD̔n 6���\O��}߾}_,� lOn�fo�      `2���;��E��J�  ��ߞ��,�9pO)�8\� �<RJ/o��gKw       �%���kr�.� l*oٱc�J���ȁ{D�`0��'���UE������J�       ����$"�^� �\RJo,ݰ^�t�F4M����� ���'N<���/���!      @�5M��xKL�C� �D�aϞ=�I)��!�1�?8�n�  `������߭�zK�      ��z�ޏG��b�7Z ��I)�qR�����`0xCDL�� ��z���\�t      �N�N�9�wD���- ��RzS醍������?�s�X� `Szq�4/(      �K]�۪��&"�/� l>9���{��O��؈��GDTU5ѿa  L�_�v��)      �C�9���]-� lN)�חnب����̼!"�Kw  �Җ������J�       �5M����� ��5H)�N鈍����%�\�՜���  6�s���7Ms��!      @9�^�))�_*� lj�ٳgϗJGl���#"RJ�)�  lj?o���N�C      ���t:���ED*� l^9�K7�T܏=����� ��������,      ����⽪�zG����- ��v����;JG�T��>�Rzs� `s�9?�i���       ƣ��n�J�  �ޛv��}[�a���{D����kJ7  DD����\�      `�><�Rz}����[  ����-����������� ��������n���C      �ѹ��#�I�;  "�3�w��H�a����I�-  �s>'�t���Ⅵ[      ��k�fD��t @DD�����4U���"�D� �������W^y�]K�       �����W��  8iy˖-�/1LS5p߷o��RJז�  ��H)�vv�������[      ���t:��9�.�lw L�w�ڵ������Akڞ� &ޣ�?�ڜs*      �_�߿_J�m��t �7���.�0lS7p?z��"�oKw  ���{��KKG       ��4����u)��-� pߘ��}W�a���{]����  �抦i^P:      X�~��xgDܯt ���ް��p�tǰM��=""����  ������X:      X�Ç��7F�O�n 8��K��T���������Kw  |���xS�����!      ���x㍋��  ���={�|�t�(L��="b0��t ���9�3�i���-      ��u��}���  ��s~u�Q�ځ����#�X� �S�WD����޽t      �z�޳RJJw  �Ɖ�[���tĨL��}����,� p���u�����!      �?�v�?�s~MD��-  ��Rz����ߕ����GD䜯.�  p?q�m�]�����t      ��v�R�݈�R� ��.0JS=p��[������  8�G?~�꺮���2      h�~����ҵ��t �|mnn���4�C����#���;  �����#      `�Z\\�p0\�]� �,^�s���#Fi������Kw  �I�y�i��\�      6��i�r]Dܻt �Y��`����6�����>"�_� `~�i���      �����������-  g�Rz������tǨM�����*  �JW�z����      �iW���fff�)� �9�C��aS܏=zMD|�t �*T9��7M���!      0�꺮���~'"_� `������;KG�æ��u��.� �Jw���v:��     �i477׏��;  ���;w�<Q:b6��="byy���R� `�έ���~���!      0M��������  k�����ۥ#�e��/��#��  kp��`�����K�      �4�v��D�/��  X�?8���6��=""�t�t ���������{�     �I�4�RJ��  k��6Лj�~�ȑ�k�)    IDATk#⋥;  ��~+++�ꪫ�Q:      &Q��{ND�FD��-  k�R����Ͽ�t�8m��{]׃�ҫJw  ��-//_�W޵t      L��i��s���d[) `:��رc�t�8m��VVV~;"N��  X����^{�����!      0	��y|D�1"��n X�+++W���M7p߿��F�5�;  ��n��w�u��t      �Y��{t������-  ��{�^z�WJG�ۦ�GD���n  ؀1??����%�G      �B��}X�����p 0�rΛr�J��sN�^��[  �+��{G��Q��r�      h�N��cUU�?"�Z� `�zϞ=?�RʥC�m������ L��󿙛�{u]כ�g:      �v�~��UU��0n &\J�o�q{�&�GDTU��ҭ�;  6��sss��9oʿ�      ���t.�G���n ؠc����S:��M;pߵk�?����  ��5MӔ�      �R������zDܫt �^XX����lځ{DDUU�J7  CJiw�4��      0n�����D�y�[  �!��[�JJ�Jk�����;  �dq�޽�KG      �8,..^���򁈸�t ����޽{T:��M���I���ٻ�/�����O�ܐLO�FQ�$�"
."����*G����u�kV/Qp����$HB2=���Cý�������g/P���\�u�W�EDP =q����\?]�I�$�������<�ӧN�W�?�  g�A��     ��;��666~;���v9��m��w��uCD�fw  �EG��(;      6�����:��oF�C�[  ΢�;���ڶ�8p�ֈxsv ��TJ��     @5Ms�����.� -Sk}ݝ��mm��#":��JDL�;  β���h�      gK�4Fć¸ h��;v\�1�#���}""ޗ� p��RzF�      ��q; �f���<x�ϳ;�����j��d7  l#w      f�q; �v�[�;��i�4��"�;�;  6C�ui~~���      ��q; ���`0�a���_���  ���;      �fyy����a� �X)e)�a����N���� ��RJ�5M���      �j����icc�7#��� �M�׫����1M���^�w��z<� `�]�4͡�      �+M�|�d2�@D|sv �f���z8ޞ�1Mܿ�d2�>"ֲ;  6�Ѧi~>;      �����y��߈�Gg�  l��Z�k�#�����XXX��R�;�;  6Y��W�F���     ����t����{J)�"� `��СC�1mܿ�Z�Rv ��R�2�$;      �?�s2�����n �
�N�U�����+�����  �;k��h��_g�      �}�Z����k#�G�[  ��o�z�?Ȏ�F�w��rMv �9'"��cǎ}Wv      �����RD<'� `�*�������Έ�%� `��WJ�OM�|[v      ��x<���zqv ���.xOvĴ2p���p="���  �*�����6Msav      �C�4/����  �b��۷o#;bZ�ߍӧO��۲;  ��C#�W_}��g�      �nM�<;"��;  ���n����if�~7�9�Z��  [�[���?p�UW= ;     �v�F�>"�%� `+�R�|����gwL3��b2�,GD��  �b߱s��_�F{�C      h��h�C���GD7� `��Z�u������XXX�xD| �  �J)7?~|gv      �p�ر��t:��-  	�7�4;b����k�  ����'O����iH      ����Gu:���Z��n Hb�|��@��4M�ǥ�Ge�  d(�\���/��      `6-..>����ND\�� ��c�~�q���2�\p?w~�F�  Yj�GF�с�      f����y�n��ø ��J)W���3t�y��PJ�9�  K)ey<?3�     ��q���kkk��n H�竫��̎��gh����k�+�  �:����yRv      ӯ�Zn����G�S�[  �����zvĬ0p�j�������  Ht��x����C      �n��x���3�  ������bv�,1p����o�s� ��=pcc�����     `:���D�|v �����ʎ�%���JD�� ��C��������     �t�����zmv ��mmm�xvĬ1p����������� �)𘍍�w�����     `:4M�k�7FD7� `
��K.���Yc�~�"b=; `
<ymm������J     �m�i�GGĻ#�~�-  S�����Jv�,2D�����""ޑ� 0%~b�޽WfG      �gqq�!�x@v �������7gG�"�{��r4"jv �4��.4M��      �����y�n��#��� �)Q;��8;bV��K�~�c��fw  L���i��     ��������ߙ� 0-J)���z��1����d���  0E:q�x<���      �ƞ={V"���  S�Xv�,3p�����sD�^v �9����G�� ;     ���4��R��� �)�[�~�w�#f���}TJi�  ��7�ر�7�=�5�!      l��i����  �6����Yg�~����j��O�;  �̣���/���!      �]ǎ���xK� |�?��z��1�|ɼ����$"��;  �M)��sss^�     h���Ňt:��DĞ� �iSJ9VJ������,ؽ{�["�/�;  ��K���E�      �w�]w�\��}_D<4� `
�277wcvD����ֺ�� 0�j�׌����      �����o����xlv �4��6���?����g��ݻ_���  �B�Z�ۖ���     ���w��q���ew  L��=��sߘ��gɁn-���  �R{'��{F�у�C      �g��y~���� �)v�E]t2;�-�ϢZk>�  _�7�R~m8��     ��9v��S#��� �)��n����&�g�`0�l����  S�����\k-�!      ܽ���Gu:�#bGv ��*�,<x���mb�~��ZG�����  �b�g�4/ˎ      �]y����xoD�?� `�ݺ���z�Yf�~�:t�"�w ��QJ���h�ew      ��VVVv�ڵ��� �iVk��ȑ#���h�M������;  �X)��aii�{�C      �b�O��6"��� 0�n�v�WgG����&����;  ���&�ɻ�     ��k��ŵ��ew  L�Z뵽^�o�;���}�t�ݫ�w ���������     �yRD4�  3���ݻ�Ɏh+�Mr���OEě�;  f����^�     ��5Msa��]�+� `ڕR�=p��g�;���}�R�F��  3�9��xv     �v���tND����u�-  3ඝ;w.gG����&�����+�  g��z�����gw      l'��2�L���n ���W�޾��7����U��� 0vN&������!      ��x<^�����  ��M&��숶3p�d������  3��k����f�      �ݱcǞWdw  ̊Z�����:���ܷ��ӧ�W� ������^�     �f�����N�ƈ�f�  ̈�w���z�0p�w^q��� ��S��     �F���{k��g�  ̊Z���Tv�v`�Ej������  ���z�i���      h��p��v�o��o�n �!�O&�qv�va�E��M��� �ҍ��.--=";     �-���^�Gv �,)��faa�/�;��-��t^��  3����W���     �Y�4�3"��� �s����(;b;1p�B�^��ַew  ̘~�ԩ7dG      ̲�x�ȈxSD�� ��:�۷����v��W� �}MӼ$;     `�F�=��wE�y�-  3掍��c�ۍ����z����;  fШi�'eG      ̚R����� �YSJy��������n��R.W� ���h���     �Y1�/�����  �A�J)G�#�#��~��"���  3补�_>q�D7;     `�---}O�u�� 0�J)W�z�OfwlG�I:��0"New  ̠'�t�M/ώ      �fKKK�L&7F��� ��RJ��]�'��z�,���  �E��K�����     �i4;o���e�  ̨c�^�o�#�+�D��WF�jv �*�����g�      L������R��� 0�j����ظ6�c;3pO4>[k�:� `F=`cc�]KKK�d�      L��h�Cqiv ��*��baa��D��&�ɨ���� ���Z�5�      ���ѣ�R��� �uӮ]�^����'���� �YUk}�h4���     �L+++�w������ �YUk}�������ܧ�m��vmD��� �YUJ��رcߕ�     �emm����� ��g��v�/eG`�>������� �v�N�s������C      �Z�4?���  �q�����ܧ�޽{��3� `�=bcc��      [iyy�Q�� ���~���������ؿ��xYv ��{�x<�(;     `+���mll�-"�d�  ̸KK)5;��g�>EN�<����Xv �,�������;      6����rD|gv ����`0xv������Z�+�  ���Z덋��{�C      6�x<~fD<?� `�u:�˲�b�Sf~~�=��  3�[���Jv     �f����Z_�� �����>��3p�N��  Z�9M��tv     ��4w�Z9"�� 0�j)��|9�)4~+"~3� ��o��۲#      Ζ�{�^O��  h����fG��ܧT��95� `��Eĉ�px��     ��j<?��:�� �����2�)��������� �x������     ��b4=������ ��J)o���W��[__?��  -p�i�ˎ      �7��a���ֈ��� �8�Ȏ��O�����G��  -P"�������     �{jnn�pD�Pv @K,���[�#�k�S���\�ew  ���"���pGv     ��ZZZ���fw  �A��3���ǲ;�{�S���}�ֺ�� ����gϞ_��      8�����L&7F��� �6(�>�����L&���tv @�R.��O��      �j&��#�a�  -��{��.;����},,,��R^�� ��Z�/---=0;     �4M��Z���  h�Rʡ�������3p����#�gw  ��7M&��     ������#b)� �-j����������ψ}��m�Zgw  ��3���#      ���p�cccㆈ؛� �����#8s�3d~~��#��  mQk}����ò;      ��޽{/��'dw  ���^��#8s�3��2�� �������_:q�D7;     �i���Z/��  h��#���3�3���,"~)� �E�t�M7y�
     H5��D��"bgv @[�R���M��3�3���\ZJ��� ��(���i����      ��N�����  h�Z�gN�>����=g�>�z��''��rv @�쬵�����9�!     ���4��Z��� �&�N���Bv�����:��s�F�_ew  �E)�Q��įv    �-����u�(�-  -�񹹹�fGp��Ϩ�.��dD�<� �e^4�$;     �j�emm����-  mRJ9������;�3�.x]D�qv @��Z�F�у�C     ��[ZZz~D�hv @��Z?���ߛ���g�>���۷QJ9�� �2.�ώ      �mii���c�  -S��� ;����}����_�����  h��F?�     ��p8�1�Ln���� �6�������Av���{L&����dw  �I)����ew      �gϞ�"�_fw  ���˲#���[�СC�o���� ��ٻ����Zk�     ��رc�YJ�$� ���7eGp���D�۽���w�  -�䥥�fG      �0wu:�_����-  mRk������������z���.ew  �M������ó;     ��777�҈��� ��)�\r���/dwpv��H�ӹ2"<�  pv�M&���Cߝ    �{m<?."�;  Z�/���7eGp��H��;G�;  ڦ��}sssew      �i8�bD��n h�:�L^�o߾�����o��~8� �mJ)G�;�-�     �왛�{YD<&� ��n8t��ogGpv��Ӌ"b=; �Mj��v:�7�8q���     ̎�x������  h����#8��[h~~���Z_�� �BO���_�     ̆���ݵַD��� �z����_fGp���T�۽,">�� �6��+���#�;     �鷶�6���� �B�s׮]��l����z[Jfw  �M���Z�O�8��n     �ױcǾ+"��  mTJ����wdw�9�[����MD|,� ���p�-��$;     �N+++�;��["bgv @}����Zv�������۷/���� �6��+��ytv     0}���.��o��  h�����gG���[n0|$"~%� ��vG�N�8��     ��h4�����  h�k>���2p�����K)�� �B�{��7Ȏ      ��p8�UJyCD8� p�}z}}��l>�m����7�Z�;  ڨ�r����ó;     �|{��=ߞ� �F��Ç�Bv���}��t:����� ��������~]v     �kqq�[k���;  Z꣫��oɎ`k�o�^�T)e>� ��J)O�����      r��N��}}D�/� ��j����p8�ak�o#�~����� �6��^=���     l��{�� "��� �Ro����/�l����#  Z�A1Ύ      �����Cj�Wdw  ��j�۽4;��e�����gw  �Q)�Y���G�;     ���cǎ�#���  -��~*;��e�u��a��3�  mTk}�u�]7��     l��h�����;  Z��v�zUv[��}:x���K)�ew  �ԅ�N��<;     �\W]u�J)�dw  �؋8pGv[��}�:y���#�fw  �ԁ�i�;;     �<;w�l"��;  Z��`0xv9ܷ��p8��D�Fv @u#�Ǐߙ     �}���"�g�;  Zj�����#�cྍ���R���  h���z뭃�     ��ZZZ:���(�-  -��^������os���E�?  �������Gew      gO��e�� ���o'O�t�y�3p��Vk��q  �����_]ku�     Z`<?�����  h�I��y�p8\�!��;1??����� �6*�|�4���      ��pة�^;�[  Z�5�^���#�g�NDDt�ݗD���  mTJ5M��     ��777����  -��ӧO_��t0p'""z��'"�� ��zP����     �޹��+���  h���#G>��t0p��<y�hD�iv @�R�7����     �s�v�G��Z 6A����~�m�Lw��p8\�t:Ϗ��� �B�R���p�#;     8sM�<)"~&� ���J)�/�خ���"�^�å��gw  {+�    IDAT��c������     ���y��UQ�[  Z��`0������;_����"���  mTJy����C�;     ��nϞ=#��  -���'O^���1p��\|�ş.�\�� �R�u��&;     �{����R�/dw  �U)�%��������;_����#���;  Z�'���fG      w��zuD�ew  �ԍ�~�}�L'w���p8���� �6���zeeewv     �嚦yZD<#� ��n�t:�����;wi~~���R���  h�o9}�� ;     �bw�Y��  h��z��'�#�^�ܭ����"� �MPk�tyy���     ��v�w\���  h��^p��/s�ܹ[���@  l�s��ׯˎ      �����#J)��  -5)��h߾}�!L7w��~�c��}�  mTJyz�4?��     DL&��#�~�  -��~��{�L?w�H��}ID���  h�奥�s�#     `;k���� ����������w�H���DD\�� �R�L&�;    �$���~�dw  �؋>���f��;g��ɓMD|4� ��7Msav     lGsss�"⛳;  Z���`���f��;gl8��R~."Ng�  ��9��     �����C#�Pv @K�͎;^��l1p������qv @K���h��     ��t��&"�dw  ����/�����w�]�vk��� �F��W���     �;v��"b_v @K��~�Cv����{���wD��E�$� ���}�޽�ˎ     ����N�sMD�� �����>��R�C�=��+������  h�Z�W^y僲;     ����ݻ?"�� �RG<����&w�]�v-D�-�  -��ݻw�#     ������Z/��  h��r�\���2p�^;p������gw  �Q�����;�;     ��v��uyD|mv @�u:��۷o�Fv��������/"ޞ� �B�R���     �6M�<�ֺ?� ��J)W�z�?��`��s6���Ύ  h�'���gfG     @��R�#bgv @�����bv�����l0|�����  h�Z��p8<7�     ڠi���>5� ��&����õ�f��;gE�߿!"ޛ� �B�����#     `�---��� �6��^���'��v0p�Y__qD�fw  �M)eaii雲;     `��Z{�� ����=�ܗeG��5����zIv @��ZϝL&���     �Y5�\k=�� �Bu2��袋Nf���U��v���� ���i�     3��8/; ���t�СdG�.�U��p����܈�=� �e:�dG     ��i���J)?�� �Bu���Av�c��Y�����R��  -����G�#     `��Z��#� �mJ)/:r���;hw6����bD�av @��Z��Ǐ���     �Y0����#�  -��~��������M1�#�yq:� �e�uuu�y�     0��a�ֺ�� �B�ݱc��#h/w6�`0�hD\�� �6���ѣG�&�     �ٞ={����  h�R�/���Ogw�^�l��'O�����  mRJ��;v��     �i���tN)���  -��~��+����;�j8��R��g�  ���M�\�     �h2��G���  -󩵵�gG�~�l��`�?j��gw  ���J)WfG     ���F��Av @��Z/��K�&���3pgK�v�m��� �6����h4zBv     L�R�+#bov @˼i~~�W�#�����p����܈8�� �"��2����     �M�<:"��� �2�<}�t?;�����-�����4� �e��4͏eG     ��X���  -R;��s�9���w��ɓ'������  h�R�����wfw     @��h�C�� ��9����Svۋ�;[j8Nj�ω��� �����՟ˎ     �,��RJ9�� �2���q(;������~��O{��>�&� �E���<�5��Og�     �V;���CD��  h�I��y�����e�����N�^���Z�'+  Ξo��    `�;j��� �6)���z�gw�=����R���s#�s�-  mQJ9t�W>(�     �����s#�۲;  Z�㥔K�#ؾ�I���>Yk�gw  ���w��u(;     �����9qiv @�L"⹽^�Tvۗ�;�����TJ��� �90��ώ     �����qqD<4� �E���dG�������\�� �����fG     �f[^^�)e�� ���?9y��˳;���t�TD�8� �-j��qyy�Q�     ��666�D��;  Zb�����px{v�3���#�W�;  Z����qyv     l���Ň�R^�� ���+����w��#���  -���x���     �����j��fw  �����]������1>���  h�Rk�";     ζ�x�Ȉ���  -q{��y����Og��?0pg��w�Rސ� �?�4�S�#     �l���2"vdw  �A)e����(��)w��d2yID|<� �%�����     8����ED<3� �%�����ώ�/e��ԙ�������LDx� �{���ҏgG     ��0�L���]  �Z�gv����RJ�n�/e��T��z��gw  �A����p�V     fZ�4O����  h�N��܋/������3�N�<yeD|(� ��w�ޟȎ     ����zEv @K����7;;Sk8NJ)?��n �u�֗��    ��j��)�����  h�O�s�9��pwܙj�~��Rʁ� �xĞ={~:;     �R�K�  Z�t�����.��dv�w�^�߿���� �YWJy�p8ܕ�     �D�4?\k�W�  �����^�������3N�>��)� `�]877���     ����  �����^xa��g����p���/Dĳ"b#� `�]����;;     ��x<���=�  3��֟޷o�&3����1>RJ9�� 0�ο�;��     _M���Z/��  h����#�Lu���x����]�v=-"�� 0�J)�{����}�C��[     ஜw�yό���  ���z������pO���L��N�Yq2� `�}������     �+��Sk}iv ���e}}�@v�S�̜^���R� � `��Z�\w�us�     ��ٳg_D<6� `�Mj�?s�ȑ�e��=e��L����#��  ����u�N�zav     |�'Nt#��;  fܕ���ʎ�{���Y����Tv �;����7;     ��[n��'K)���  �aݻw���po�3���g'��s"�f�  ̨�ر�@v     ��'Ntk��ew  ̰�666~j�����C��2pg�:t���k�;  fU�����r^v     DD�|��ϊ�o��  �U�փ������������� 0�������     8q�D7"�dw  ̪Z�;���_�����;3o8�^J��X�n �Q�뮻n.;    ����o��� �+�������gw��`�N+���?+�\�� 0�t�ԩ��     l_���� �[�'��O�z������� g�>��?|�S���"��-  3�O�ӯ{��߿�    ��s�y�=3"^�� 0����OdG���;�r�9�0"�4� `}�d2ynv     �S���v ���������:U]Y*pw� �>�F�#���b �Y��Ą- �@C�:�{���+KHwWUk�3y0����G7��AŇ���"�MY�>tU׹��s#f饪>gy>��ׯ�s��u���^o5;���;e߾}�N��'">�� 0������ʎ     `�����@D|Gv ��hD<��R�C`+�3q���j�K�  c��ʎ     `��� �k��h���C`��3�����J)���  C��m;�    �t8t�Г"�q�  㦔�����dw�v0pgbu:�gG��;  �I��a���7dw     0fff^��  0nj�o���n���b���Z\\�l�ӹ."ֳ[  �I)�Gڶ���     `�>|������  '��O�����ٳ���������v�Qk��� �1��w�S�#     �l���n  3���<{������T�`��Z�����#�� �qQk}�cǾ�m�av     �gee�j�o��  3�5Ms ;��ܙx��:77�����% ��TJy��ݻ���     `2�×d7  ��w�޽�ǲ#`'�3>��t����� �qQk}I۶�     �R����.�\�� 0F>{��ݻ�;�X����v����  #�:??iv     �e8�n  '���4Msgv�w��`0����  㢔�#�     L��~sD\�� 0.J)k�~�u���ܙ*m�gggo���g�  ���\^^���     L����~ث  ��w=ztv�4L��n���qcD�� �1�c    �3v�С���ސ� 0&���{ڶ�Bv�4w�R�4o���dw  ��K:���     ��N�Ӎ���;  �A�u����ߟ�ܙZ��-��  c��Rz�     ���n��A�� �qPk���~��; ��;Sk�޽�����Z?�� 0�J)�9r��     ��]�v�0"�� 0�lff�%tL5w�����?�E�fv �������fG     0~ڶ=����� �1�Z�U�n���!���������RJ��� �QWJy����Wew     0^�;�gG��fw  ��aD����?���!"����K)���  e��s�?���     ��w�1��  c��MӼ!;F��;DD)������� p?J)�<�;�    ���}hOD|cv ��{�����fG��0p�{8p�3����|v �������fG     0J)Mv �������u{�����Qa�_dii��J)�F ���n۶s�     ����Ջj��:� `�m���>�����D�׻="�Kv �������#     m��pv �(��v���~?�F��;܋�`�/"ޙ� 0��m���     �^-//?&"�� 0�~���*;F�A
܋�m?��t�����[  FQ)����fw     0���  ��������0���>t�ݿ*�<#"jv �(*�t�     =�������;  F� "�ZXX�;;F��;܏^����֕� �������fG     0ZJ)7E�lv ��zA�4������c��Zߚ� 0����Bv     �cmm��Z��  �����4��ew��3p�ж�]�v=5">�� 0���v�mˎ     `4?~|oD<(� `��ѣG��0��$�t�M/�\�-  #f�����#     �׶�l���1 �?�陙��ڶ]��q`�'����A��G�;  F�޵���#     �5??�����O �j�/..�Mv�w8M�,�Z�[v ��9}}���     r�R~8� `��i��ʎ�qb����R����� �sS۶��     �X]]�w��� �QRk���`pkv�w8E���?��t�Dı� ��ݻw?%;    ����n  1���xF۶��7�p���j�O���� 0*j���     v����7E�%�  #dPk���[n�Tv�#w8M�~�u��۲;  F�cVVV�    ���ݰA �G����~����W>.�=z����  ��C     ����ꗗR��� 0B^���^�����@۶ù���k���n ��+:��     ��p����  ����=��0���-,,�]J�&"�f�  ��������     �����Y�� ���'N<uϞ=��!0��a4M��֧G�0�  [����n��A�     l�����"�k�;  F��N�s��7�|WvLw�"�~����� ��{vv�Y�     l�}�  #��Rn�v����Ia�[��뵵���� 0^ض��    �	u�С�dw  �������28�-TJ����ƈ�O, `�}������     l�N��� �l�����gw��1p�-�������"��-  �J)7     &���Wew  ${����3۶f���1p�m����WD\��-  ��t�ȑGfG     ��:��"bWv @��gff�r��7ߕ����I�4�mv @�������     �����Y����  H4��^�������Tz��+"�� �,��g���~yv     [�����G��dw  $��~���0��a�R�9��xwv @�Z빵�gew     �e^�  ����^�����t�����7����,"�>�  C��Ew�q�Lv     g�СC�SJytv @�Z�{w����RJ�n�Ig�;`qq�o"����LN ����×fG     pf:�΋�  �|fff�򅅅��C`��i��M����  �Pku�    0�VWW�."���  H0�����_e���0p��4͡���� �O\]]���     N�p8|AD���  �i���MӼ!����;�RJ�t:ώ�?�n �ae8�0;    �S���vVD�Pv @����z��0m�a�u���onn^�n �aO�+_�e�     ���Ǐ__�� ��J)o���id�	�����R�eq,� `��ڵ�Y�     ��d  찿�״m�������z�?��gD�0� `���Z�#     89����-�<:� `�t:����Od���2p�DM��J)���  �A߸�����     N�p8|~v ��R��v����if�ɺ���#��;  vJ)�a    �x�+_�e��=�  ;���z�������R�`0���x{v ������͎     ���ڵ�ٵ�s�;  v�O7Ms$;0p��ж�fgg�RJ�Pv �����ynv     ���Z"�y�  ;����`��;�P������ʣj���e�  l��ݽ{����ݻ�    �?�����xcv ������w.,,|2;�np��������Ԉ��n �f�b0\�    ��+�<?� `�]k�ܸF��;��^������ ��Vku8    0�VVV.��^�� ��6k�����wg� ���;���in����� �͞������     �S���E�lv �6[������s�0�v����Z�[�;  ��=�$     ���o�}WD<;� `��T�4�!;�w�0���ݻ���quD| � `��Z�y�����     ��`0�*"�� ��~w0<?;�o�0�n��OE��qWv �6yPD\�    �?��^ �$�눸�m�����Èk��/:��u��� �J)��     �8r��#K)ߛ� �M��t:�7M���!��3p�1��v�XJY��  �&�:|��Ɏ     �v���Ϗ��� �ND�5�n�=�!�3p�1���Vk��gw  l�R�s�     �����9��� ��PJYh��M���1p�1r�ر����  [�����n��A�     �j8gw  l�Z�r�������3p�1Ҷ�����U��� ��Tk=wvv���    �i�M `B��c��gG ��������ݝN璈�Hv �ۛ     0������Z��;  ���g�m;�N��;��n����pxED�[  �пZ]]}lv�e`    IDAT    ��)�썈�� ��>Xk���m?��:wSKKK�3"�Dĉ� ��2=�    �����Ϊ�>-� `}jss��~��������k����dw  l������ώ     �����D�Wfw  l��Rʵ���vp��a������Z��;  ��y?�    0-j�^� &E-�<����vvpf�a4M�TJ��� ��Pk}~v    �4XYY��R��fw  l�Z�^������3p�	PJ�G�}N)���[  ���:���#     &�p8|nD�� �-������`k�Äh��Ǐ�""�Wv ���t:��    �Fm�ΕR��� p�j�o^
�	b��[n�������� �3����Ύ     �T���WF�Wgw  ��wonn^׶��`��ÄY\\��N�sY)�s�-  g�N��';    `R�R��	 ����R.��������;L�n���Z�3#b�� p��     l�Ç�ˈ��� �3p��rI���pv���aB5M�˵֛�;  ��w���<*;    `�t:��� 0�6"��^����!������.��*� �<;;     `��q�3�֧gw  ����iޔlw�p\p�M���gw  ��Z��������     �w�y�E��� ��Qk}Y�4�)��^�0���ٳy����#��-  ��ˏ?~Ev    ��1;  �4�R�4/Ɏ ���;L��m?733seDܙ� p�     l�����*�\�� p~g0<��R�C��g�Sbqq�o;�Υ��� �SQJ�pee��    �q���������  8E���ظ�m���`g���v�冀^ǲ[  N�LD<#;    `<3;  �}��rɁ>��w�2�~��J)�Eĉ� ��Uk}N��dw     ������Dģ�;  N��"��^����`g����z�ώ��� p���#G�7;    `\�Zo�n  8Y��ϕR.o��}�-��3p�)�4�ϕR~4� �d�C�/     ��m۳�y� `l���{��d� 9�a��z�WD�Ofw  ��k����ώ     7���WEėew  ��ZJy^��}v�����`0�F�k�;  N�������    �qSJ�B& 0j�z��Oew ��aʵm;O��7e�  ��0     �`yy���}�  '������#�|�@�m�>77wMD�iv �xܑ#G�    0.j�7�} 0���`0xQv0|� ���p���ܓ#�/�[  ����泲     �A���R��� � ~{nn�m��C��`��o��G�ǳ[  ��3o���]�     �nyy�����  ��]333W-,,�F��;�O,--} ".��Av �}�������    �1���  �����p������f� ����g����Z��_q �H�.    ��;|��|)��� �������/--�]v0z܁{����7F�0� �^\q뭷~Ev    ���t:�F�y�  _���Z�����v0�܁��4��SJY��  �ssss�fG     ��Z�3�  ��F)��~����`t����뽺ֺ�� p/��     0�n��EĿ��  �5"���vߘ�6w�5M��%� �K<����ߜ    0jv�����	 FO�i��Ɏ F����R��ݻ�o�n �b�N��    �QSk�& 0jV��YɎ ƃ�;pR��ݻ1�)��-� ��R�Ѷ��    �{���|WDx� %?�������0NZ۶���ظ���?�[  �������͎     no F�?TJ��!��0pN��7�|׮]�.���e�  DD�R�     DD۶s�'� �o�����m��!�x1pN����'777/��;�[  "bϫ_���#     ��޽������ ����s�9�)ǳC��c������d8^�� L��>���_�    0�x	 ��wnll\�o߾Av0�܁Ӷ������'G�g�[ ����    �j��z�W�Z/��  ��_��'8p��8m������,�\�m d�����͎     �277w}D�ew  S�#333.--�]v0�܁3���������8�� L�������     Yj���n  �W���q�����d� �����~�ͥ��G�fv 0��     S�ȑ#�,�<:� �Z���>�i��e� ����2�^ﵥ�gGD�n �ҷ���<*;    `��8q�� `:�R>7/_ZZ���`r�[����lD�pv 0�j�q    ��Rk-����  ��F�������e� ����rM����xiv 0�n��;f�#     v���꿉����  ��f)��MӼ!;�<���h��%��� L���y�ߓ    �S�l	 $�����z���L&w`��z�~)����  �K)�a    0ڶ���k�; ��RJY������ &��;�mJ)��.���n �ʞ���s�#     ������#⫳; ����^���L6w`[�ٳgs0<-"ސ� L������     �͋� �{u�4/Ɏ &��;��ڶ]הRޖ� L�:    �D;|��|D\�� L�Z�����`:�;�m�ϭ��_�� L�K�9���    ����t��ew  S�W�;vc۶��`:�;��������0"ޓ� L��O�8quv    �v�^� v�o���]߶��`z�;jaaᓵ�﫵�7� �l��;    �DZ[[��R��gw  �̓��ʅ����!�t1pv\������̅�� `����>4;    `����_�� ��*��~��ʶm���Lw E���h)�	��� `bufgg�ˎ     �^� ���O�8qq��?�L'w M���pD<!"��n &S��!    0Q:���� `b����ƥ���?�L/w U�4w��#�c�- �D��Ç[v    �V�t:7DD��  &ҟmll<��������;�nii�/#��Z�'�[ ��t]v     �zjv  0��?;;{�q;0
܁��4�_D��Għ�[ ��RJ��Z�ی    ��w�Сo��o��  &�_���<ᦛn�xv@��;0B���;����Għ�[ ����+++�Ύ     8S�N��� �V�3".\\\����d������?��^G�[ ����    ��f  �õ�'4Msgv�3pFN����R�E1�n &��m��    [+++�ߐ� L����'���f� |)`$�z�?���#�Xv 0r��~wv    ��R% �U>OZZZ�@v��1pFV�4�O��/d�  ���8�    �R۶�Z�� �D��Z��������b����i���t�ǳ[ ��Vk�Ӷ�lv    ������ވ��� `�}6".������?����v�o���`Dld�  㫔�U�{��ew     ��R�*�3uw��yr�4��@܁����_�Gĉ� `|u:�@    �X��eʫ�; ��UJ�\D\��vߑ�p2܁��4�/�R��� `l]���vVv    �ɺ�eʯ��  �ֱ�pxi�4��p�܁����~6"�G�[ �������'gG     ��N�s]v 0��_k}\������Sa����i~9"�n ��S�     N�=/R>%� ?��7�Z����3��T�c�i������n �K���Ç�gw     <��Ǐ_��  �ί;v�)�~�Xv��0p���������>1"ޟ� �����4;    ��t:�=� �����શm��p�܁�v�M7}|ff梈��� `|�R���     pVWWϩ�^�� ��R��:���m۞�n8���[\\��N����lv 06.Y[[;?;    �lnn^�ew  c�=�N��n�����3e�L�n�����."6�[ ��p������     ����\��  ��Ow:�+]
Lw`b4M�[�fw  㡔rmv    ��Y[[;���� �X،��u�ݿ��*��D��z���;�; ��Wk�xmm���    �/u���'E��/�TJYj��� [���(��z�9�<'"�2� yg���_�    p/��  �¯w��#� [���8���D���� ��Rʵ�     _���o�UJ�,� m��u:�g�Rjv�V3p&R�4\JyEv 0�j����y�    ������ `�m����C ���;0��=��Z�[�; ��v����/Ɏ     �G�֫� ��Vk��~������b�L��m��N���� `t�R��n     ��h�v6".��  FW)�m��W�; ���;0�z�އK){�; ��v������     �{��E�Wfw  #�Z����ٳ���܁����^[k��� `d�}���K�#     :���� �H{Q�4wfG l7w`*�u�Y�"�� �h*�\��     L�;�c&"���  FS)�uM��\v�N0p�����ݵ����� ��K����ώ     �ׇ?���G�Wgw  #��Rʋ�# v��;05���["��; ��t����/Ɏ     ��p8�:� Y�n������b�L����ň�Dv 0zJ)�f7     өm�N)��� `$�n��{Mv�N2p��-����fw  #��Ç�gG     ���������� ��9>33��K)5;`'�S�i�_��_��  F�9�N��    `��ë� ��SJy����{�; v��;0�N�8�dw  ���zUv    0]j�%"���  Fλ�;�C� f� 2���o��IOz�"���- �Hy����#��;�s";    �����]JY��  Fʰ�z����! ��L��`���� `��7??av    0=:���� ����~�o�L-w`j�m;�t:{#b#� ����    ��Pk-�7I �+�|�s�����L��T�v��*��fw  #���o�}Wv    0������  Fʋ���7Ȏ �d�L���>����� `d|�ѣG�    L�R��� �Hys������l���۷oߠ�rsv 0:j��    ��pUv  026"�E� ��� "���/�Rޖ� ��Rʕw�q�Lv    0�����#"�!� �֟l��}� ��� "J)5"~8"6�[ ���5�Ї�;;    �\�/I ��㛛�/ώ � ���zZJ��� `dx    �6�V�A QJ���o�+�`T�|��Ǐ��Oew  #��ZkɎ     &���ʣ"⛳; ���'G�����Qb��En��OE�˲; ����#G�<&;    �<����� `$k��ڶf� �w�/1^���  �y"    �&�d  �J)?����(�`��|��mO�Zo��  ��Z��n     &����R�� ��kff�G�# F��;�����o��_��  �}������    L�R�S� ����7�t�ǳ# F��;�}��6��  �p8�"�    ���˳ �t�۽{���# F��;�}���,��dv ���j�    l��>$"�� �*��߻w�Fv��2p��N綈�Tv ����+++dw     �ovv���(� @�?�v���0�������gK)�fw  �JDx2    8c^� ��aSJ�� ����=z�U��  �C'    �L����O��  R������gG �:w�ж�zD�$� H��#G�<8;    _Ǐ�$"�; �4�333/Ύ � '����bD�Iv �f������    ��*�x) ��kߛ0�NB)��R�� @*�O    �i����wE�E� @�c333/͎ � '����v)����  �\���vVv    0~��'Dă�; �4+����0.�N�p8�G�0� H�{}}���    ���t:^��)Uk�����Jv�81p8�~����_��  r�ZB    ���Z"��  G���񅅅��; Ɖ�;�)*��8"��� �R��F    ��#G�|GD\�� ���G��&;`�����iWgw  )������    `|�C/C��*��ܶ�zv��1p8���Ogw  ;���0
    8�g  )���v9;`���|�ֺ�� �Rʕ�    �x8r��#"�_ew  )^\J�� ������E�'�# ���+++ߔ    ���pxUv ��J)��4͛�; ƕ�;�i������ ө�zYv    0�j�Wd7  )~4; `�������WE�ǲ; ��UJq(    ܯ[o��+"�q� ����^���� ����t����Zgw  ;����?�?�5�    ��:묳.���� `gu:�g7 �;w�3t�ر���  vTgss���    `t�Z�	 ��M�n��� �����m��R�m� ��r8    ܗ���s"��� `g�×e7 Lw�-p����D��; �u��Ç�#    ��Sk�0"�~ S����KKKo�� �� [�m���p�; L�sJ)n`    �/@���������Ia��Ev������� ��rH    �m�v"�� `G�j��}Gv��0p�"{��ݨ��<� �Q��m;�    ����;�q�� ���a3�������🍈�gw  ;�+�9�    ���Z��`���i�?Ύ �$� [hϞ=�����)�
    �b��˳ �SK)/͎ �4� [��ѣ����  vF)��    `4,//KD|Sv �c���z�0i��X۶�Z�[�`z<����ߖ    �����F������;�6h����� `g�R��n����{{����;�]{�$���<I �@[�c�ql��#!m���_Нk�����ԧ��f�S\�pHB�8$�@��!�$���<q�� %�Ȓlyf�Ջ��H������{�^��r�>{-    Z�?e  #��C�});`�A)�F�]� �h�Z�cv    ��رc?o��  F����;�# &��;��\v�eG�; ��+�\s���gw     yz��[� ������Ɏ �T����{��"��� `$J��sv    ��-� �h���۳ &��;�mݺ���; ��px    Sjiii[D�lv 0���?�0���h���gJ)G�; �����i��    �������+� �N���v�!3p�~�o���dw  C�c�Ν7eG     �Wk��# L��8p�� ���`����Nu:�_��  F�!    L�Z뛳 ���ϥ��0��F`yyy)"���  ��?d     �u���+#�� ��}��ɓʎ �� #����݈x{v 0t�9r��    `tz�ޯd7  #q{�4���i`�0"��c���� ��9�   �)��tޒ�  ��O�<��� ���`D������ ��,    ���~���Z���  ���rg�4�ew Lw�ZYYY���d����n{Av    0|333o���� `��YJ����ib�0B�~���[� �Pu�n���    ��u:/:�������}&�`���X�׻="V�; ��r�    �����Z�/fw  C��^�����ic�0b���_��dw  C��i<K    ����>"^�� կ.,,|7;`��$���5� ��o߾���    `xJ)���  �3[�n}[v�42pH077�W��?��  ����%�    �Z�d7  C���������id�����ݝ�  O���    &ԑ#G.��+�; Ŀ+�    IDAT����nw);`Z�$�������|v 04�^\\���    `(�Cv  0<���8p��� ��� ��  ��-�    0�|��	�����n �f� �v���ވx"� �\    0awD�M� �p�Z�r~~����if��h߾}�qOv 0����瞝�    ���R~>"��� G��9�� 0���-//�'�; ���v���͎     �ˍ 0���駟�`v��3pHv뭷~���� �pt:�]    0!j�%"ޜ� ͯ6M��0��Z�����������    �1w�رk"��� �P�XYYqI%@���������  ����Ύ     6����F �P��������� ��d1;  �N��+�    �����Z��z����g������x(� 
�^    0�_�dw  Cq|aa��� �?w�v�;;  �7�u�]?�    lʿ; �T�� ����EN�<������ `�:��7gG     ��t�� ��C��Ev ?`��"M��#�ײ; ��p�    c�i���֟��  ��zwv g3ph��'O�+"��� V)�����ew     �}��=�+� ���:u��# 8��;@�4Ms:"ޞ� ��3g�ܘ    �_����� `(�6M�ώ �l� -����; ��*�8   ���� L��<y�# 8��;@������� `�j����     �����OFĿ��  �MӜΎ �\� -���ߖ�  V)姎;���    `]ޒ  \����� Vg��Rsss�� V�����    `]ޜ  ������>;����X)�׳ ��s    c�i��u:�=� �`���{� 8?w�۲e��Fķ�; ���٥��m�    ���ܹ�Z��� `�=}��'�# 8?w�ۿ��R���  j�����    ��x� &�ۚ��gG p~� -������X��  ���P    ƃoy 0YN����+;�3ph�����#�#� �@9   ��[\\�Ɉ��� ���Zkaa�� \��;�(��-� �+�9ryv    p~�N痳 ���v��5���3p�/"�:� �R�/e7     �Wk�# L��fgg�o ƀ�;�����  `��   @K---m����; ��)�ܓ� ������'O�'"��� F���wH    �̳�>{SD���  �ɝ;w~$;��1pMӜ.��;� �gΜ�>;    8W���# L�Rʯ�۷o9���1p#�^�m���  �!    �P�շ; ��u���Ȏ `��������"�� �`�R�   @�,..�dD�2� ���r�-�̎ `���L)�m� ��\y�ȑ˳#    �p1 L�Z�=� ���;������È��� ``~1;     8��; L�R�#sss��� `}��L)�F�۳; ��qX    -����-"n��  �ײ X?w�1��v�YJ9�� ��6M�5;    �x���]D���  ⩧�~�xv �g�0�8�T���� �@�ڵk���    @Dxq &F)�=MӸ@`���~���� `0j��    �|����� l��;�����8"��� �C3    Hv�ر�Eī�; �������������Z�od7  ��;���    �f�~�E 0!J)��n `������̻J)��; ���v����     Ӭ�j� ��镕��gG �q� c���O�Z?� ؼN���    �4M�5"n��  �w>�tv g�0�:��'� `�Z�{�h    ���ر��E��� `����-��3ps������~9� ش];v����    �R^X�������G�# �w�	��t~3� ؼR�C4    ��� L��g �y� �̙33� ��9D   ����_ZJ��� `�Nmݺ��� l��;�x�[��O�� ����;�,;    �I��-� �@�o���'�# �<w�	QJyGv �y333���     Ӥ��K� ���Z#���0p�����fw  �f�    #r���n���� `��znn�ϲ# w�	QJ�~�
 �ֺ��Z�;    `<��WGďdw  ����  ��`�lٲ�]��� lB)�_;v��    ���=� ��=��t~';��1p� ��r�7#��� ���z���    `��}�� `��Z?0;;��; w�	���=� �oOv     L��ifJ)7dw  �SJ���0� fnn�#�k� �ƕR�4M��5    �ݻw�>"vgw  ��>��`L L�RJ-��3� ؔ�ر���    0�z���� �����R�# ,w�	����ΈX��  6���p    ���rSv �)˵��ʎ `��&��Ç���~2� �8�k    0<M��D�� ��||nn�[� ��;��zwv  �q�֛���?    ��]����; �MyOv  �a,0�N�:��Tv �a�߾}�k�#    `����� �M��֭[?��p�L��i�-��?� ظRʞ�    �D�NgOv �)�ۿ��� ���`��z�wg7  WJq�    ؽ�޻��z}v �q���d7 0<� l~~���Jv �a7?~��    ���ɓo��� ��=z�С�dG 0<� ���;� ��]��c�]�    �ˉ 0��]J�� ��;���ޓL�� `c:���6    �Z�� `�j��e� ��`�:t�"�� `��d    ��h�fkD\�� lا����>;��2p���wg7  v���ǻ�    0	�o�~mD���  6����� ���`
����G��� `C.}�'�Ύ    �I��v�d7  �L���Pv �g�0���N�Z� � ؘ^�wsv    L�Z�� `�>������ ���`z�;;  ذ=�    0��E�u� ������d7 0� S�ԩS_��  ֯�r��޻%�    ����ʛ"�� `C�|��^��� F��`J4M�/��vv �!�N�8���    g��=� ����޽{{� ���;�tyWD�� `C�d    �83p����t\�0E������."�<� ؐ=�    0���y^D�)� ؐ�����uv �c�0eJ)��n  ֯�rý�޻%�    �Ѯ]�����ew  �Wk}Ov �e�0e�{�ߋ�3� ���<q���#    `�Z�d7  ��e˖�eG 0Z� S��[o�ND|4� ؐ=�    0�J)7g7  �?o��ofG 0Z� S��M 0��   ��=z��Z�Ogw  �WJ��� F��`
�޽���O� ���R�o�fkv    ��Z��DĶ� `�N�R>����L�}��-�R>�� �O�u����ߘ�    �ֺ'� ؐ���>����L��e  ���tn�n    �qRJ�M �P�ն`J�L������G�7�; �uۓ     ���ѣ��Z�� ��m۶�Qv 9���޽{{��dw  �SJ��i���    0z�޵�{ ���߿�Lv 9����� `��Z��޽�u�    0J)7d7  ����mZ ���;�;x����� ���Z�   ���� ��ۧO���� ��L�RJ���?� X7�r    pǏ�Fě�; ������i��� ��L�n��I' 3��k�%�    ���_��k#��� `}lY 0p�r���_��  ��w�u׿͎    �6��z	 ��?��%/y(;�\� DD��+ ��n�{cv    ���; ��R��������  ��; ��vߛ�  ���9    ����  ��%� �q���/G��dw  �b�    �q�ر�G�K�; ��+�<>;;��� ����� ��+��ΟȎ    �6���.� �1Sk��RJ��  ��; ���7� X�����    ���`���}�3� |�����"�s� ��8�   �U�� ������Ɏ ����Z�_����ޘ�     ms�ȑ�R^�� �]���� ���; ���t~/"jv �f���;.͎    ���!"Jv �v�nץ� |��; �w�����R�4� X����̛�#    �Mj��g7  ��7���_̎ �=�8K��/b`�ܐ     mRJ�1� X[ �b��Y����#��� ���;    |�ѣG/����; ������ ��������#"���  ��ڦi�fG    @�Z�����(�<2??��� ����s�R>��  ��%�v�z}v    ��`��ZmT 8��; ��v���^v �6�~���    h	w /� �}�8�-���͈��� `mJ)�    �zǏ��Z���  ��K���� ������Y 74M��;    ��c�=vUD\�� �M���� �� �*�| "jv �&�߹s竲#     ��`�t:���n ���X����^k�\v �f�    �j� 0V����|v �d���|(;  X3�w    L�� ����~��R�; h'w Ϋ���� `�n�    �,w�u�+"�'�; �5s�" �e��y���5"�&� X���}��/͎    ��n� 0>�q�ԩ�fG �^� \P���� ����}O0   0�j������`�4�� ������$ ��R��    �ķ1 ����n ������������ew  k�f    �Α#G^���  �䩝;w>�@��pQ��g7  k��cǎ�Hv    �R��ƈ(� ���Z?�o߾�� �����*���x�����Ɏ    �Q*�\��  ��G� h?w .��.{8"��� \\��a    �ƥ 0�۶m�ǳ# h?w .j�޽���� ���);     Feiii[D\�� ��}���?�@���&��g7  krm�43�    0
���WG��; �5�Hv  ����59u��'J)��; ��ڱk׮+�#    `���`<�R�G�# � �I�4�k����  �ġ    S���[ ��G<��� ƃ�; kVk�pv pq�V�z    L�� `<|$; ��a��z|4"z� �E9�   `�;v��#��� ��J).U`��X����oE�g�; ��z�ѣG��    ô��� ���ggg�*���a��z�E- �_���Ύ    �a�t:�f7  Wk�h)�fw 0>�X��e  ����^   �D��^��  ��G� /� �ˡC��_��  .��b�   ��j�f&"���  .��ɓ'?��x1p`�J)��  \ԵM���   ���}���FĎ� �>�4ͳ� �c ֭��?� ����K/����    0�n��� `MlL X7w �mff澈8�� \X��w�   �D��^��  \����ǳ ?� ������Dğdw  �   �	�r h�/,,,<���1p`�<! ��   ��s�m�� "^�� \X��c� �'w 6���},"jv pAW.--�Ύ    �Aڶm�uQ�; ��ry" b���>|�Ɉ�Bv pA����7fG    � �Z��n  .��^~����x2p`3<% ����     �� ����Ͻ{���; O� lX)�SR �r�Vw    &F�4���j! ��M	 f���=������  ί�zm��dw    � �޽�ʈ؝� \Poyy���# _� lX�4���	 �X)�_;v��    0�^ϋ� �~�ַ����# _� l�'� ���:�   `"�R|����%`S�ؔ~������ ���   0A|���+���)� l����7"�� �9�   `�;v�G"�U� �=���O�yv ����M��[ h��wdG    �f�z�k�� ��MӬdG 0���� �@�͔R�Ɏ    ��(�x� �φ�M3p`�v���PD���  .��    c��zmv pa+++�� ��3p`���۷�gw  ��   ��Uk-� �ݗώ `��0(���v�.;     6���~eD<?� � � �������av pA?~�ȑ˳#    `#J)o�n  .����0p` ����>"��� ��C@    �U���� ����t:dG 0��R�_�@��   0�������}&;��`����Z?��  �_����    `���y^D�:� ��Of 09��n�{D��; �ՕR^�4�Lv    �ǎ;���-� ����1p``8�TD|.� X]�u��;���    ��(��!� ���.��G�# �� �'� ��ޘ     �tMv  p~��������� `r�0P�VON@�9   `ܸ� ��V��2p`��m��pD<�� ��s�    ��{�ggD�2� 8����Of7 0Y����������; ��jiii[v    ��3�<����fw  ����Ç���d1p`�j�����ں����    X/@��qv  ������v�� �b�~ߡ     c���[ ��� g����8q⑈�vv p^�d    ��@��z��� �<� \�4�Z맳; ��zcv     \�w�qiD��� `u��/>|��� &��; C��t<A �u�ѣG/Ɏ    �ٲe�"�dw  �uv  �����p�; ��L��{]v    \H��Cv p~�N�6��0p`(<���fv ��R��A    Z�7, h����� �L� E)�F�� ��j�   h;߰ ���r���'�# �L� M)�ST �Rn�   �͎9�xYv ��Z��� L.w ���rv p^����;weG    �j:�� ��\z�0�04�RD|+� XU���^�    ����� �b�N�� &��; CSJ�� h�7f    �jJ)� �^������� &��; CUk�$ ��5�    ��Z��; ���� L6w ����  �   �:w�u׏Eċ�; �ՕR\v�P�0T��bD|+� Xտ>z���#    �_*��1� 8����� �l� U)��Z��  VUz���#    ��\�  ���/,,<��d3p`��  ��a!    m�w h��� �|� ���� ��J)o�n    �����A h�R��; Cg���:t���� `Un�   �5���"�ǲ; �խ��ܟ� ��3p`�J)5"��  Vu���⋲#     "bffƋ� �^_=|��� L>w F�U �^��k�     "��b� �e��H�0�V�� @K94   �-j��U@K�~ 0*� �ġC��6"���  ���   �6����x}v ��Zk�?;��`��(}:;  X�Og    �����#�� ���<??��� ���; #�* h����;";   ����v�4 �e����02�n�?; �R333   HUk}}v p^�g 0=�����GK)�gw  ��:;    ��� �Sw F������~:� 8W��u�    L��� �U���C�����0p`�j��e7  �2p    �ѣG_/��  Ve��H�0R�^�S� ��.����4;   �����\�  -�2C F����ZXXx<"��  �Qfff<   @�R��� ���+++dG 0]����� �B   H�� h��u뭷~';��b�@w h�)�Z    IDAT'��    dq� �P�����3p`�z�ާ� �U�.;    �鳴��;"^�� �����0r� ���Ç���G�; �s\�4��#    �.�>��UQ�; �s�lٲ�� ���; )J)~� �e���WdG    0]:�����>���� Lw R�Z����ݮ�D    F�7) h'� R������5� 8�U�    L��� �s��}w R������_��  ��0   �����{�D�� �9�K)gG 0��HSk�K_ h�Z�U�֒�   �t8y���-� 8�g���NeG 0��H��t��}v/..�<;   ��qUv  ���� �^� ��v�DD��  ���v_��    �Ը:;  8W��0���e�@�[n���hv p�~���,    F��� h�^���lv ����l~� -SJqk    CWk-� h�R������2p U)��� �n�   `�9���� �l�V�����le  �xɑ#G^�   ��s� ���
�f�@���]D�cv p�Z��E    ���� ���ʊ�; ��HWk��� �l�N��"    �� �ϣ�~2;��f�@:O[@���   �as�; ��C� `�@�N��`v p��    �m����Z�e� �9\R@:w ҝ8q���tv p�W5M�=;   �ɴm�6, @�z=�����tMӬD�g�; ��tw��yev    ���j� �������ˎ  w Z���+ h���    �L� �>��K)5� �h�N��+ h���    �L�w h���  ������������ �,   ����m��� �l�w Z���V���;���  �rU�4�o   `�VVV^[�; �(��>q�� �`� @��%0 �ˎK.���dG    0Yz���� ��j��i��� �0p�]��efff^��    �d)�\��  ��f��0p�5j�ED��  ��   ��*��6� 8��; �a�@k���}+"��� �@����    L�Z�� �Yz�^�3� ���h��v1p   ``�=��x~v p��>|��� �g� �J��� ��eKKK��#    ��~߅
 �2��� �_2p�U��u�����    L�R�k� ���Z�n ����V����jD�cv ��V�j   0�5@�t�]w Z���֩��iv p��    �oM �._=p���hw ���  �,   ش�i:�����  ���v Z����)���	 ��5�    ���۷��ֺ=� ��Z�f7 �3p�uv�����x&� ��-..�(;   ����t\�  ����  �a� �ξ}��K)�dw  gyuv     c�7& h��/���/fG �3p��j���n  ���   ���	 ��/����ˎ �f�@+�R<� -��t>��c�~���{����'��!�"*�\�Z�o�1������z�C�F>�-���^�K�J1�����샤1Ɯ�}H�������
�O���]   �=���c�i1>�$)�0UQ 0!   ������Lv ��0U
� Lҋ/���R�f�  n��Zkd�    `5moo?[J��� ��l6Sp`���2) �����O��dv    V�7�  ���Ǐ� �D��)Sp�	���    |^�  ������ �w ��a
 &���   ���� L�0F�,w &�ҥK?,�̳s  7y�   ��r� 2�͌0Y
� LV���K)�g�  n�	   ��}���=ZJy2; p�Ս��ײC �N���Z�/�`:���~#;    �ecc����� ���^x�jv ؉�; ���� �遭��g�C    �Zj�� bl��Sp`���C L�|>�Fv    V��; L��A &M��I�ַ��f)�w�9 ��"���    X9
� 0!��:w &-"j)�g�  ���    �I�U� ��ӧO�2; ܍�; �~� �1   ��������x4; p���  �Qp`��`R�>s�̑�    ���0�  Ӣ���)�0y�/��!; PJ)���g�C    �2�`Z�%;  �F���;q�ąRʛ�9 ��"��    X]�)��t�k�?� �Qp`U�� &b��gg    `5�Z�`:^?y���! `7
� ���  \g�   �e�Z���?�s  ��Z���X	�08d�tX�   `W/���S����9 ��"¸  +A���p�ر�K)��s  ��R�8{��#�!    ���|��� �Qp`%(���{�E��G�9 ��a�ki    �*"��� ��/��Fv X��; +#"~�� ����     L��; LǏ"�f� �e(��J,��t(�   �wH 0FX%
� ��a� `:<N   ���f  n2*��Pp`e�<y�祔�9 �R��K   p��������pv �:�� �w VFD�Rʿe�  J)�;{���    L�0�  ���K/�t>; ,K��U�b ��n�X<�   �i���  LDD��ƨ  �w VJ��G� ���p   �wG 0� �w V��; LG�uV�    ؉�; L�� +E���r��ɷK)��� �Rk�jv    &�8 LD���� `/�X)QK)�7; PJ�H	   ���?x���Dv ��Rʇ/���;�! `/�XE�,�i�j��Ε    ���W�>[J�� ��v V�" ��G� �RJ)������   ����� 0����Qp`��f3�/ ��Z��    �wF 0FX9
� ��'N����6; `�   �;Rp��X,FX9
� ������ @)�֯fg    `Zj�F `>8u�Ի�! `��XU~� +   ������x:; PJ)�z; +I��U�� ��w�    �t�С�K)��9 �R�n +J���4��}e ��o��_�   �4�f3����w V��; +���ӿ,��&; P��Ɔw    ���" �� �*w V�/�`"£%    ��] L���N��uv �<�XY�V_�4x�   �}-;  PJ)��d ��K��Uf� &��;    ��jv  ���Щ `e)����ap�iPp   �|���}����� (e�fg ��K���u�ԩwK)�e�  �S}��   @�����eg  ������� �y)����  �졇z&;    ��� ��?O�8a0�����J��*���Z=^   �� �A������J��gg  J)/   �Wk�Zv ��R�k� �^(��҆ap(�iPp   � L�. +M���v��ɷK)�s  /   Z��+�<TJy<; PJ�u?��  �B������zv �<���3&   @��������� �O>��㷳C ��P> `�E�/� Y����>���    䨵�� L�k}��! �^(���j��eg  J)�x�   h�0�#; PJ)��e �{���:Pp�	��>��   ��n &����� p��Xy�.]z��2�� ������    @w ���Pp`�)������RJy3; �΂;   @Ӟ�  �ťK�~� ; k�� �ς;   @�^~���J)e�  �O���� ; k���Zv �<�ꫯ�   ����?��D�� kA���0�w �w��ŋOf�    `\�� �`�u���Z�w ����<f   4fwB 0�X
� ���'O����~v h]���   � `677-���X�V_"@2��   h�;! ����?�Av ��X�� �<f   4���tv ��L �6�X�V���|~G   А�_~��R�Vv h�Q@ ։�; kcccC� �=���Fv    �q��5��iЙ `m(��6�x�7#�rv h܁���'�C    0��l�~ 0��܂; kC�����s�-j���� Z�X,<j   4b� ����>��g�! �~Qp`��" �E�GM   �FD�� ��z��Cv �_�X7�e  ��;   @#� �$`�(��V�aPp�d�V�]    ���>�� 0�zQp`�9r�R��n@.�]    x��+�le� ��E�w ֊�; k����R���9 �qO�}��   ��u��5C �o8x��g� ��I����gg ��mnmm=�   ��5�͞��  �_����������� �l{{�z   ���� $�	 ֎�; k�뺟dg ��u]�q   `�E�;  HVkՑ `�(��v|� ��q   `�E�3� �u
� �#w �Α#G�,�\�� ��	   ��j�Ogg  �@ ֎�; k����.���� g�   `��9s�K���� и�<�Fv ���XW�P�\u�ܹYv    �G���  ߛ/����� p�)���~�  ���;�<�   ��1��� ��? ֒�; ��! �E�_gg    `��� ��`-)����ap��|V�    ֔q �� �%w ���˗�*�|�� �   `ME�q H6���������Z��~(��4; 4N�   `M�Z���  ����SO�<; �w �V�կ�  �/   �5��+�<ZJ��� ���s�=�� �A��u�W\ �멾�;   ��իW�*; P^�  �E� ���u�w ���C=���!    ����;�� Z�� �3w �����w H6�Ϗeg    ����>�� Zg��u����:u�ԯJ)�s @�f���N   ���� �u]g������ڊ�ZJ��� вZ��    �_q,; 4������� �E����X�D;   �O�Ղ; ���� ���Xk�֟dg ��Yp   X/}�w��'�s @�����Xk� �5/   �5r�С�K)d� ���`�)���f���; ��ʹs�f�!    �?f�ٱ� к�Pp`�)��֎?�A����9 �a�~��'�C    p��c $3���Sp`��r rmnnz�   X�z  �G'N�x/; �'w �^D�r �p,;    �ͱ�  вZ��� `�)���j�� Q�ժ   ��8�  ��� �~Sp`��Z�� Zǲ3    p�3 �\: �=w ֞�; 䪵��    ����~����9 �e: �@�����o}��R��s @�����   ��9�R�Fv h�0
� �=w Z�Fv  hU���W_}�@v    �! ���S�~� ���; ��3 �]�|�+�!    �g
� �("ވ��� ���; ��� ������    ܛ�8�� g��&(��
�< �e�   `����\� 4A��V8�@"�^    �� ��} �	
� 4��ѣo�R��s @�j�ǲ3    poj�� QD(��w �����o�R��� ����'   �
���`)���9 �a����� 0w Z�Kf Hb�   `�:t�/�� d�E��W�C �>h��; �y���    +h6���  ��y �
� 4#"���  ��G�>�   ����  �8w ���@K�  �b�8��   ��'"�eg ���< �w ��u�� $��fV�    VT��� ��y �
� 4�ĉJ)�g� ���ev     >7w ȥ�@3�h� $��   ���� @�߽��Kf� ��(��w �s,;     {w�̙#��?�� ���  0&w �Rk}#; 4��   �jr� �"B���(�Д��U3 ���ٳge�    `o��{2; 4���h��; M��f�j�<1���";    {���  вa���w �r���_F��� Ъ��
   �b�ap� �j��h��; M��~����� Z�u�w   ��t  ��cǎ�� cRp�E�l�<־    V�; ���s�=�� cRp�9��7�3 @�j�־    V�; ȣ� @s�h�w ��1   `�D�; Hb��)�М�l��� �0��   X!�����Xk=�� Z�u�� �Qp�9׮]�Yv h��/   ����a�  �Z�h��; �9}���Rʇ�9 �Q_����   ���w H4��; �Qp�U� ���ѣV�   V��; ��t����C ���h�ϲ @��aPp   X�. ��,"jv ��; M����3 @��~   ��a�� @��I
� 4i� ���   �JQp�$��@��h�l6s�$�Vw   �a�  R�6 �$w �t��U� ���   �
��F)�� ЪZ��; MRp�I����R�G�9 �QV�    V�?��?>ZJ9�� Z5�͌��$w Z�Kg �a�   `D�{ �������� �h�/� �#gΜ9�   �])�@��GD� �hV�Ղ; $���    �]��/�3 @�t h��; ͊���3 @ì   L\D���$�� 4K��f9@�_    ��p  ��> ���@��� RY�   �>w8 ���:�} 4K��f���K�R~�� Zd�   `�j�
� ��h �Rp�i�V���~o   0m}�w��ǳs @�"��'~�� �(�д��K/ �a�   `¶��+�lf� ��Zߊ��� �(�дZ�_z@�    �X,�� @c} 4M���E�[� �Q���?x0;    ;�> �c���)�д���3 $�t���    ؑ�; $�7z Z��@ӆap(�$~s   0Q�Vw7 ���:] ���@�N�<��R��� �(+`    �n  ��; MSp C Ha   `�"�� ���'��gv Ȥ� ��";  �H�   `�j��gg �F���~� ��h^��|v hQ�u_��    ���� @ Pp��u��� ТZ�gg    �O}����B)�Pv h����<w p8�a   `� @��8�� �)��<�����/�Z#;    l>�+�@��0�@��h^�u�(��� Р��|�;�d�    �O�� $Qp w (�w�Y)�7�9 �E�X
   01a� �\�rE���)��u� @����R   ��qg 9>�����e� �l
� p�/� A�u�   �ǝ �8�  �@� �;�  �   `z,�@�| P���RJD���  -��*�   LL�U� r(�@Qp�RJ)���! D��R   ��qg 9j��3 �(�@)e6����  -��   0-}�,�|!; 4�8 w (��r���wJ)Cv h��]   L��֖A ȣ� E� J)����WK)�e� ��D�S   �	���	  �b�x'; L��; ��3 @�>{���    \
� ��ӧO_� S�� 7��W_ � "��    �M�� 9t �w ���; ����)   �tXp�
� p��; �Pk=�� Z4�GS   ���w5 �@g �@� ���� ���:�    QkuW 	"Bg nPp�666�gg �y4   �� �F� nPp�>��R�"; 4H�   `"j�
� �`6����  S�� 7<���ۥ�w�s @�<�   L@��])��� Рz���w�C �T(��-j��3 @�,�   L��Ç�TJ��� ��������  WIDAT�! `*���� � �    0����  �:�  �D� nQk��/ �c7~   @�Z��� �Q�
 p �ED��� t��|$;   @�"�  �� �B� �د� @����x
   �� ��U �[(��sh��0|9;    � ��U �[(��-��C# $��k   �|�0����
 pw �ũS�>)�|�� ZSk�   �� ��A� n�� �� Ƨ�   ��K� �Aۗ/_�Mv �w �M�U� F�eg    ��������� �D� n�u��; ��ϲ    ��W^y��r4; 4HG n�� ������ ZSk}4;   @��� ȡ� �Qp���Z`|P   ��s �CG n�� �� ��    Q�u�g  AD��< �F� n3��; ����3g�d�    h�?�@ ���; ���>sx�V�    ��Z�� @ ���; ܦ��˥���s @kj�V�    ���Vw ���; �ٻ� �AQ   �D�w ߕ_|�w�! `j���|! #��#*   @�Z�� ߯"�f� ��Qp�;Sp��Yp   ��n Ƨ�  w�� w�fg �yD   H�`|
� p
� pg� 0>w   �$�Vw �n ܁�; ܙC$ ��J   @��ﻈx$; 4H7 �@� � ""`|�   lnn>\J�e� ��DĻ� `���>���wK)5; �dw   ������ 	����)���}���av hIDxH   �ax  (���)����s��q=r��9��   ��; ���'N\� S�� ;����� ���|8;   @���  ���  0U
� �3w �l6{4;   @�,���t `
� �� 0���m��    #�� 0>� ؁�; ��:�I YD(�   �lw2 0���I �(��,�����   �ϝ �O' v�� ;p����    F�� )t `
� ���b�0	 �Sp   �; ��= ؙ�; ��ʕ+�Rjv h��T   �����f3w ؁�; ���k����s @Kj�~�   0�3g����� ��z�꯳3 �T)��ݽ�  c-   `D `|WO�>}!; L��; ܝ_���"B�   `D�V�1 0��"�f� ��Rp��Sp�qY   �0�c `|� p
� pw� 0�#gϞ=�   �!�`d�~v �2w ��Z��; ��o�   �Sk�bv hM���� `���.��Sp��E��3    4�] �,"t �.��.,����ax8;   @+��s ��E ��Pp����� Ff�   `<�0�������Sp������� �Q   `$a� Ffl �N� ��ԩS��R.e� ��X   �����677��.�`wV�`DU   �Sk�� �_�p��! `��`��i Q�u+;   @C� ��>��~� S�� ���*���"�j   �x�� ��t `w
� �;�K QDX   ����z��r$; ��_�`w
� �_O��j�
�    #�z��{ YD��� �N� v�u�� �1V   F����pv hM�U v�� ���� �1
�    #�A� FVk�A �](��.f���% �K�   `� F: �w ��b�p��qm�}�
   ��j��`d�`w
 ��Ç;\�����   �Sp��u]��  �Pp�]|�߼TJ�,; ���
   �φa�Bv h�|>Wp�](��r>�  -�����
   ��"� ���>�? �](��"�� 0"��    �/"�E �u���k�! `��`	�Vw ��;   �������q� ��`	
� 0.w   �QXp�q� ��`	�	 #�A�   `�)���t `	
� �� 0:w   ��� Fd\ ��� Kp��qE��U   ��g� Fd\ ��� Kp���)�   �Zk�R��s @K���r�`	]�9d��,�   ���>ZJ�e� �����(����C& �hw   �}t�ڵ��3 @k���r�`	p��Yp   �_�0(��Ȇa�= �%(���?~����� ��   �� ����; ,A� ����av h�1   ���� Fv��� X��; ,ϗ� 0���Ν�e�    XW]�meg ��|����� �
�`y
� 0�x뭷�   ��j�
� 0.� X��; ,�a F����`v   �u�^ `\: �$w X��& ���:��    ����� FTk�9 �%)���"�a F�X,<�   �� 0�� ��Pp��}�  Z�   `�Xp�qu]�s  KRp�%���� Вa<�   �Z��� ВZ�� ,I� ��u݅� ��    ��� �N� ��� K�� ��l   ���� �� X��; ,�a ��   `��Z�fg �����)����a��� Z��   ��ܽ ��j�: �$w X���}M �:�    `�)������9 �%)���^xᅫ��ϲs @C�   ������f���; ,I� �Ɓ FRk��
   �Ν;7���� -�x� ,I� ��Bv  h��;   �>x��,�Dv hȕ��d� �U�� {����Xp   �����] `\� �
� ��V�N IDxh   �����] `\� �
� �7� 0�    �`6��w��[< 썂; �ͅ�  ��    ���z4; ����`o�`o:`<
�    ���:�. 0�Z�1= �w ��N ��V   �}0�{ QD��=Pp�=p��Q��޹   �>�w �� 쁢  ��0� 0�x��Gg�    XCG� @Kj�� �
� ��`\���G�3    �� 0.] �w ؃Z�� Вk׮yl   ���
 ���`o�`��s���f3w   ����z4; �d�X� �(��<xС F�X,�   �Z�; �w �w ؃��ۿ������ Z�u��V   ��,"ܹ ������� V��; �AD�R�'�9 �[   ����  В�����j�r�X� wT�=�����>�%�1,�"q	��
�IHȆ�{2����/R5�}'�]+3��� ���= ��e   �)ܹ @��߿�  A� I�wO (b�;   �� �����p�= �� �� P���   `<w. PGc  Iw ���� �("���    ^��� ��h  I� I��� P$"^͞   ���  Dc  Iw H�;|@�;   �x�\ ��� �$p�$�; ���&   0�� ��J< �	� Ͽ����V   ��>~��� �2�5� $9�@ޏ� ����   0�ϟ?ݷ @!� O� I˲8|@�   �\.w ��1 �$�; ��| �{p   �z��o�Z H�@R�ݿ��HD��   0���� j��=  �� �� P'"<�   ���� �e�; $	� iY�; i���   0PkM� �,��<�; $E�W@���   t>�� P�= ��@Rk�� �xp   �z�Z(  �,��$�; $]�W�; ��   `,��V�]c  Iw H���u��"�w�    ��ܷ @!_��<�; $����| Ա�   `�eY� PKc  Iw Hz���O���� ����
   0�/�@���� I� �8�@���{�   ���< (����/ �$�; l?f�  �߿��
   0��� �Hg�  {#p�z�̞ ��r��   ƹ�  �����:{ ��; l#p�"��Y�   0�� ��k�  �Gw ؠ��
 E�e��
   0H��w �cy l p��eq�"���]   �w- P��< �@� �� u"�w   �q� P��< �@� ��B���|��
   0�� P��< �F� D�C( �^�6�   �Zs� E�E� [��mlp�"6�   �c�; �i�� vI� �����b    ���HD�g�  {$p�m~�  �����   `����� `�� ��� P�w   �A, �R�8 `�; l6�@��p�   0�M� P�� `�; l�{�� ���γg    xAܵ @��� �	�`�; �qv   g�=  ȫ>��= �H  �i� ���[�    �q� ��9{  ��; l��3 �Q�   �r� ��u�@�� 6轿�= Ekͣ+   �8�� �Hz�w H��!p�"6�   � 
	� O� ۼ�=  ��   `(w- P("�1{ ��; l�Z�@�֚GW   �q�� ���� Iw � "�:{ 8�eY<�   �� �Z6�@��+ l#p�:ή    �X&  ���  �F$  ���Hk�<{   �D� �� �$p�m��  �""�    �k�Z��  �F� ��� E�    C�k�Z��>}���! `O� �������tz={ 8�޻GW   �qܵ @���Ƿ�g �=�@җ/_�~�
 ez�~w   �� �XD�6{ ��  $-���3 ��D��W   ��~��Ξ Jg  	w H��Ϟ �D�   0Ʒo�ܳ �: H�@��' �{x   ����= ̡3 ��; $�� �<�   �Z[g�  �3 ��; �9x@���   pss� &�H r� ���	 �z�^   X��= ̡3 ��; �9x@-�    ����3 �A�  A� I���� �Hlp   ����= �q7{  ��; $-�b�	 ��    ��g�, 0�� ��@R�]� �\�   �� ��Z ��@��_ (��   `�eYܳ ��d 9w H��0 ��   `�; ̱,�� � ��Zs� ���   `{, ��k� ���
 y~?��K_   �1�����~8�N���������#�!�� ��˵��?��n    IEND�B`�PK
     ���Z$�3  3  /   images/7ade412b-fa94-47ea-987a-d6c9baa14438.png�PNG

   IHDR   d   �   {��n   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��]�Uy�f���o�'YB�D��[��Z,� B���c�6E%�S�֧�$��XJ��Q�Z�h}
�<-�#�XD�b�f�Mv�ww��ߙ���3sw���͝9s�ݻ��/{�ܙ3��|�9�s���"��{�,W�\�r�J���[�%�2����,���"Kv���=�����F��t�X�gYǲ�����%΢��X��fy��,a�S�w!�ES�c����.I��Pﰏ��{Y�ay��Y^f�W�W@���K,og���d���_����%I��$���4�����7^����;�2K4x����7n
�1e���d|��f
z�-7��X^a��X�c����D�����3Kd؉DXַ�Ί֌���;X�IV�Hj��,��Ĝ��E:�p,�SD�Q�?G�ߨ}��BѠ�L�rEc-���s��ɸ�,+c�Ҥ����Z,
�5�_��cq�-��i\M�3l��>��Y�H��W��繐���!����(+���NQOG��QT�Ε/�\8����l�Q*&'bl���#�C��̘��g��#�� CC>A2,���d��1����"��%���Y� y�% �шF���ζ�l<�4U���<��_�9�岘�%�#`�*cj�f�}�U��S B\ځ�6�oPiq��^��J	u��{��ՃS~4��@��n�.&�0eu#k0M%��|�D9!K�(�q��5*�"3?ux@Kt�c-�%��~��2ۙ����d͈�d���E�5+���<2��)�9@>�f�X2���Y��D_���:���s4&�
�~2K������ P%��T�e��JG!�� ��5�N]�C�'���͋�'�C����E8/ЄW�)�+��!{5�Q���l�K�͖Q�[�&(Td9������;���yd8@c���k�:�J��>49+���t$��,��H��.��k�� v,H�T�ĩ����F�S�!�y��`�����&e'S�����}�(�د;!'xh5y�X�Z�E��PL'�b��?�B����W`u?VC1p�ɣ�Q�[a �e#/Q��CsB��/�۩ق�`��P����O����k�Q�΁DX���g�E1d\3�E�a�;��+�iё�zӰ!`��F+� Yy��$�p�����鲿x���Me� �`B�|����|�~�򘘩�u%E�9�C\h�k�i*:�p����h<B �eӵ��1Jƣ�4em�O��)�ȭ�lhb� �I��6ߛ��u�Đ��!d��@�������4;����!�Ў<��hV�&���E�o�v�źh�"�/��ά�Z���iJ���E�/�\伣Nh�0W�Y��U�"�@�Y��\�E�/Xl��g��!~`/�����i0��(G�f��1�ri��b�R�o��XX]O��-RO��"���DZ&�a &���ݢE�_訲�İA�4�%ur���ei�%��zb�@���U���r��t�LH�<q��]�dZb/�4[EZ@MD��]1L��J]�R�h��K���N�����7!֬FZ���*Z�@�h��Y�8��_��}b���>>�כ�t6[�Y�l�B��;z�EP��-[�;_@����}������hk>� ���I>�W��-ш�#H�Jщ�b6��du�%��Yv�-Wp�#�9/tXb��q_REK�zXC�wdŦ;hb�gjN5��l`IA3��(���!�͞�V���)t��銑�`��a�!��u�=y�H��J㿤�u!G�w��,�C7�y,#���~A	A�8�a)�Q]h�k�GE��|��tir�B�����.��{,y>�����&\u���$9�y�@l��4]�i�����]�!.s�M���G�wٰ�PGk$��(�Q"���vZ�R��zL���?���gĊu�GGZ��&&R0�J����R9/�Ē2M-�wş�|��kJ.��\O��x�J�#��D�S���l�@��I�ɫi��7�z,���C-�&̍�oT�a���)��� B"���I�&B\ځ���T|��#�TyK%�JFPs��
3�����n!{z+?í��Iu�Ι��|X���<��M���!�	�۴��w��1S:&!���G���$�Gz;��8� 6<#ܑ�;l��'@��
q��cg���1;A:�n�J��̊���}�خ ��k,�{�X�4��I�>?i�[ly������3y��Q1���4kE�u�Yʑ���$��Z\��5E �ɇ'�)�k�[-Z�(!�ЬL�Qn,�m�ܲv�A���_���y\��fnRF����:�^2X�Hv���.cy���x}��|AB*��N�����31/�ݡ���6B41�1�S���RS"m}�cڠ�XbeJ�d�:��ɚ�V&$���4� !��A��{�A�Tl�������"(��T�&��Q���8�D8�Gw��z�
Ŵ,A�$�R:��@D�m-6�J��T��ibT���I�]b��3�"�?2][^a�
�#Æ���"�����@
̗	�e��K�`��_�u��d!2>�r=*?��ۓWvS")�*]��*��C�cT��3rrh�hd8�df�.!L��,=х>
�I���>=�>I�����
B<d��e���̝��+��] d z�L©{��	���?7�" >bB�.�@E��F��,�,n4���rY��a s���h�*�T���w�B}�~�%�z^;�%���@T�}cS�i��2���oNx��1�����f�(,-I��C���$�~��t���~����D��P�㝎�=L�_�?�qoR&ģ�Y�S���S��̹�-�^����{k���g��烀�	CD�}.��d�k-q-���̖��lt�b6}y�<��#���J�.��F�¹	���` 1����4��aqf5A�>2��4�C\7�3tp"#*�6.4�-f#��1�ׅ�j���	����S�¿a��$'pWV\ �S�cV�x6]F9$�����q?��������hb��s��:��d���=����!��wy��7�+@����\��=$=�(�9N>��?�e����a9Я�Ͻ��Xu�h�WCnd9O�֍�µ2@@&_���7��$�|a��vT���
�^"�����4��$�-��h����x���&*��W�&P"����c�w�o�v������Y|��(�b�7��6Z�,���b{Y%�OY~�D��{)��E�U�A&ٟa����H׊�+*40)�"�Jk��k_gM�O<�qkȵ,g:_�@��;9��t&��G��n�ʛ�$ىN�ѨA�L��a:� 1'^�7����7�0c�3|��}��f���O��k�{�?��ڂ�l���^A�:4{·��D=1��݃[��Mz�,�x�\*F�O�^/���	�Wj� �↪q޵�)� %��^�D̿�w�޶��t�!/ź�}�t�Д*w3����0,�X�a���g�j�6g�D���ϟ�s���Y"Ok�'-σ`n�WF?W8^�q�C�5Ւ�]ۀ1Q�.r����F��!3��^��6˃��6�����k��o�lZ�A���WX"0�x���h��#٣�E�]��+�\NUa?U˥�j�Ŕ��D�wn-�K�$`��Ti��L-
����ihX(��P	�\��-\#�}i���Xb�pX�)���d��$�@:�3Q���9��v0x�b�Q�qL�����x���}�G���.Ie�,���L�	b4Y�̑!֐��"�:\N�5I����B.7�h��Q�@�yLB[����4�2�2�3n�8��d�)S�ӑ�I#i�F��-��~���/ɏK�s��Ig���7���׼	��E��i4����Q�[���e��!O�M:��pt��a�vVt��ͼeU��6�P�h���������J������"��@��r&�"�X�0��Sn2xHAO#i	�(ru%u:wu��<�>&"j�\�loG�ϟ���������W8����o���K�v�Uq���ʎj�3B�uE���������E�%�����-�5�D��JR�Yo�`��D�����bI��c���\��sڞ���7�})+�7��֚!������t������'^�S�dM2)7ιB$lxH�sN��F&��DT��xF��\�Y����Y8�(Y��T�d
�[�7S�4�tњ�s�}��i������F�g��ȣ�nWˋ3냿|j�]���V"�`-sq*:u�\*h*l�>~i��93�go�nn2��#L�Eo;9���^��$�o��(��z�^1o?|�B�B�S����dr�f��"L6�n}�B��y�
�A�>�YVd8@�W�s���W!�L����9j��j]�!+��/ [�p�]
!�
	`�'���z뭴\q�-�Ў�l&Y'��LL�B��%�V�	�ܹA	I���o��o���͉�-A�N��Du,�҂��*�!V��7J�Iʻ;�
���f&��:0�����:��[��r�ݡ��AR�`5B�@2X�w6�Aj@]�Pp�A��E�����B�@���{/e�Y��{�!ϳ\����X>��-G��"��R�� �i��RH�͏���LˉW�`sS�b�O���Hmv	|���z�<��JhZxȀ��c�I���@��X�UH��{H����>�ҡ��<��`2�mR#��i�-�of���,Pq�; %g�"Ac����Y��|_��5�-�d1�|B��"�B�X��E�;ї4)2���!%����a� Z� �8w����@���(��k�r���Mȿ���u1��R0������\@�I48/���/Q�\�}�_A���&J_`-��M����ĥ�~����� H�B�x�~��i���n����B�J.ER<��&�_1y,�~�}@�� �bї��:`������|:����6��P��S�ǂ�]_	����Ѻ��;�\2�߷o�����!�F��}ރeB<Z�U�Kɳ�[d���U�ti����r�CL�*p���x��xH���L7���V@��4�$����nr�x���B�������\^7� ���R��]O ?R�{I�邁[���ظ�$#���_	����k'--\�rb�`���5�@�FYUC<�`J�-�����I�7i�r}i�19�p�s`!����g&�k�ϊ��5`��͖�܈�uiI"(C9��b�^4L��Lb�d�Bư(�ii yU�
������X�𘁔=�``�B��TK��+I��L-�o0~��}�����빦�������@]=�炚�8 ��I�� ����F�G\� A�TGW_v>�Z� �����U^����]jl\�x=,���5����1b�D��3�zC�C�=��~�@�W�e�B�\b_�,5&�&Q��@PBT���pǼ@�	�m�b���!.��5Dp��0�G��e�B#u�}�=���B�.[P��-,�S��O�Rc�M�ףn�U^N�,˻�_G�ռ=�BB~Lj8��y\7�	I$�ϋ}�/��v881��PcktU�ˠN^
z�oB�l��t~X�R��$p4�q�h���p��nVTLn�wz%-�m5
��ur4��*�`^��DH�0Wq��)�p=�$��>B�1��U�5���P�UB�I��xP͓R����LC%�J���'��/���"��aB5OJ��?T�
V    IEND�B`�PK
     ���Z��F�} �} /   images/b63deb06-c33f-4ae3-8f73-25229955b1c1.png�PNG

   IHDR  �  D   CzWF   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���{��y^�'�U�Y�s�����xYD�F@P��;�Ჱ�ll쮷]5aa�V$��uB�n�0ܼ��������,������Ow�S��2뒷�#+�T�S��\��WY��Dd����'�'N�y�����   @�	I~>�J   `!���3�<S:   eUK   ��OK��(�   P�S��zs�    ���  ��ޒ�g�|b�     ,�7$��$�[:   �(�  ,�?��ǒ\-    �'y_��(  �2j�   P�W%yg�V�     p�F�/O�����  �9Sp  X<_���'��    �QM�G29�����   p��  G%��M��    p�U�|v�ߐ䇒���  �<(4   ,�z��L򕥃    �#xO��%9(  ����  p��d2�ꭅs    ����$_�d�t   Ύ�;  ��v=ɏ'�=��    �)��$_����A   8
�   ��'&��I>�t    8E�$��I>\:   ��Z:    g�w'��Qn   ����$?��3J  ��)�  \>oM�I^W8    ���I�M�/(  ��U+   �S��$ߟd�t    8cK�{6�*�  �S��  py��I�i�f�     pNjI�x�^��+�  �S��  p9��Ç�   �h*I�p�V�S8   �I�  `�}K���ɉ<    XD�$oI�II�[6
   �C�  `~U���$�t    �@~ �ےJ  ��)�  ̧z�wfr�    8�}I�<�A�    <w  ��SO�I��t    ���]�/N�+�  ����  0_���7��    s�?fr,m�t   ��;  ��XI�I�R:    ̑&��$/�  �kSp  �kI~<��/    �Ї3)��z�    �:w  ���$�6��(    �سI>7�ӥ�   p��   xUoJ�3Qn   ���	I~.ɛK  ���  .�OL�I~K�     pI<��'��g��   p2w  ���S��?�o.    .�k����@�    �K�  ����I~&�[&    �o-ɏ&���A   8N�  �b�=I�M��J   �Kn5ɏ$����   p��;  ���Ln�|�t    X�$?�䏗  �D�t    �$_��2�    ��z�/O�t�_*�  `�)�  ���I�?�iQ    ���e2�]�  �0w  ���d��I�T:    ,�Z&��>��g  XX
�   �L����A    �$I5�I�J�   �(�  ���    ��;  @A
�   ��OdRn_*    8��;  @!
�   �K�    �C5ɗ$�p��  ΍�;  ��Qn   ��R�d���;  �9Qp  8_����,�    <%w  �s��  p��0�&i�    <�i���$�T8  ����  p�� �r{�t    �LK���;  ��Qp  8;��    p�Ԓ��(�  �w  ��񇓼'��    p�(�  �!w  �ӧ�    �۴��kI>X8  ����  p���   `1(�  �w  �������;��     �B�  ��)�  ��v    XLJ�   �H�  ��)�   �bSr  8%��   ���&��$��A  NK��H�ٜ���jY^^>�O�s�ھ���T���륥����{�ܥ�����Z���۫�jZ��}�W*��ۧ���~��888H��?�?ooo/���^����� {{{�֍F����[���������h4�o��`������\ �9t��O%yo�    �J�  ����$�:�z�  @9��˩�j���G�V+�J�XI��l޳=9�P}R��V�ssΓ��GK��j����џ��\F����=%��_���e0�^��^��ce�����*�O�?Z���ߟ�����?��E�n�a>6 p��%��$?Z:  �<Rp  x4�=ɿKr�p ������=e񥥥Y�{Z����l?Z@����I�z�~��>��ۛ�f�ƙv`��P�����p��x<+�-�O�G�G�?-����������t���?}�i�=  ��n�/N�S��   �w  �����L�7� �mZ�>߽<�>�P~�>�{��<�}&���~�?+�O�f������|������y�t���� � v���$?[:  �<Qp  x8o���'� �"x�ݞM,�N+�N:�N_^^N�Z��?�����d�ݯ�qMK��i�w�~��$���I�t�����i����f8foo��G��[I>/�J  �
�   �Z��'���A ��f3�Ng6�|�|t��t���������3�|� xu���t�|�׻gB}�۽g:�t�`0����=S鷷�3J< ��+I�P�_,  `(�  <�+I~*��(�ӳ���f�����,//�^���j���N'�z=KKK���v{V@o�Z���'m .�i�}ww7��`6I~0�����g?{{{������z�{�3-����Ϧ�pi��䳓|�t  ��N�  �u��D��(`ѝ4��t�N�s�4����v�=������Z�V�# �׫M��N��n�{J����l�t���݌F��`�}4�<|  �>�  ^�R���t% ´H�l6�n�ge󥥥c��ѧ�ޯ� �㙖ޏ��f��"�����b���M_�P>�I����A   .*w  ���'yO�/.༴��,//��j��jeyy9�v{�z���j���dyy9��˳������ ���������������eoo/�����z��ݝ=�ۺ��׻���}M�ȯdRr�t  ��H�  �d�$�J򕥃 <���v�=�����2��~����������Z���(  ,��t�����S�N�?i����́$��$ۥ�   \4
�   '�'I��t�r�V��I�G��O�����cէ�wOTo6��?
  \�~6!~gg�ش�����z��z�ٺ�������f8��(����I>?�^�    ��;  ���A�?_:p�M'�7��٤����O���G�]__O���  \D��(����&������l�۷og4������I�8��j   9�
  p��&��J� �G�ٜ�ϧ��z�>[wA���z��(�  �lZx?� �<t�ty{{;����G ���%y[�q�    ��;  �-�7�<������GK��v;�v;�V+�N'�Vk�  �"������nz�މ��'�O���g`��#�W�  p(�  L�wI�a�j� �hN��~wY�u  ���j��.�����F���a��I��t  ���  �?��;��J�y��%���������  �ˣ�㷶�2KǇy5��.��\:  @I
�  ����I�/I�t(�R��J����-]�n�S�8�   ���������3{L_O��G�����$_�䟕  P���  �"{K�K�)N��&�oll�ʕ+'NS_[[K�Z-  �� S�oݺ�����>������i$�ϓ�`�    %(�  ��%��$�J�W����������euuu65����N'����t\�  ��x������������v������[:6���$_��'K  8o
�  �"��$�w�7����t:���x���W�\I��.   .�n�����{��O��O�O��ߺu�td�f��N򋥃   �'w  `�\M�I>�t�_�����F666f���$��֯���R�Oq   �G�~?�nwVx������f677O\�֭���ұ�/&��$)  �8�  ,�N������j6��	�G'�}LK���   ����?�?]w�������ұ�x�N�I^.  �<8  ,�z��%���A8{G���b�݅��E�����j�ұ   f��i���+�-��z�ܾ};�Ѩtl��J�$;��   �5w  `T��;��J��4����fcc#kkkY[[��^]]=�����F�Q:2   ���F������N����������lmmekk+�oߞ��}�v���JG���D&<��   �%w  `|k���t�k6�������FVVVf��	�G_����R�OX   ��5���v���9�����N677s�������&��$��A   Ίv   p���$�t�E�l6��t�n�����+W�̊�W�\I�ݞٯ^��Z�V:2    ����+��z�ܺukV��.�z�ܾ};�Ѩt�E������!   Ί�;  p��Iޙ�Z:ȼZ^^���F���f����r�ʕ���fuu5���Y__O��,   ���A�������۷oϞ777�������ܾ};�o����N���o$���!   ΂�;  pY�5ɏ&Y.��»r�J��ַfuu5W�\��766��   8�2�t:���Vnݺ�_��_ȇ?������(�W%���A   N[�t   �3𻒼'���>��e_�e�c    �@��z�\��+W�[�h4�L5�?K�B�[8  ����   p�>1�'Y/d^����
   ��acc�t�y�L��I~G�    �I�  �L6��X�7�2O���JG    �$�U=��$�:�'�  pj� �ˢ��I~k� ��T,    .
Ǫ�SI~<ɕ�A   NC�t   �SPI�]I�`� �h}}�t ���V��T*��\�TR���y�I�ﻟ�h��x|���px��x��x<{߫= p~�zd���G��5�~�(   �G�  ��^��(b^��3 pT�VK�ZM�Z�-�j��.O���'��_��>��%��`��h��h��p��p8[�ߺ�2  fuu5�jՅ����g2�O%���O  �9��  ̻�1�_(b���3 \~���G�ZM�ј-���4�T*��q/�ii��l>������>2^u��I�  ��R�duu5�o�.e^}y�oJ��J  xT
�  �<�#I�n���m�`~-�O��G�^O�V�MV��J�2�o������-�������������� �e������x�J������A   �3  ��zs��I�hc4I�4��Z��1 �����~R����A����I��� `^mll��h���[�|4ɏ�  ��� �y�T��&Y+d�mll��  �R�+�7���s��L�Z-��V��V�eyy������X���� ���988H���x<>��  �OE#ɻ���$�_�,   E�  �7KI�e��P:�e��� 8k����>}LK�J�tD.�J�2���ݦ�����Y�}�|ppP - �q
�f#���|F��g  x`
�  �<�d2u���rY8Y ���4����,--��lfyy�$v.��*�O��O'�O�M} ΋cV�ꓓ�H��N�W8  �Qp  ��7'���!.'����>-�O���̻J�2���Q�� �yr�����$ߙ�O�  � � �y�g����!.����� �B�V�Y^^���R���g˕J�t48W�+��F�Y�}oo/{{{����h4*� ��:_���I�f�    �E�  ����%�$;eN��Z�X�}yy9�fS�^E�ZM��J�՚��{����^vww3& �cVg�o$y&�;J  x5
�  �E�[�|O�f� ���� ,�Z��V�u���h4JǂK�~��fޕ��W���^:�eUI��|8�O�  p_
�  �Ev%�%�Z:�e���"�T*i6�i�Zi��Y^^��x��f��f��u��� �^/������x<.� �(VWWS�V3�JG���I~ �g%���Y   N��  \T�$?��SJ��VWWKG �SW�׳���v�=��^�VK�NP�׳��6��r<g?�^/{{{��� �b�T*YYY���V�(��F��%��$��  pw  ���I>�t�����w�j�X���j�V���<�J�����,//������fwwwV|7� .���U���30�9I\Q  \(
�  �E��$�t�ˮZ�fee�t x(�B{��J��I��2�.�z������݇F�Q�������n����݌F��)�Ӷ����{�t����%��$_Y:  �Q
�  �E�UI�z�����(p�U���d�v��v��J�R:PP�Z��}p�ڵ����������eww7��tL �1������(ޖ�W�|C�   3
�  �E�$ߖD��8I�ET��f��v����%�v�UU*�,//gyyyVx���K��Sx�9��չ��$O'yg�    ��;  pq��$�I�*dQ8I�EP�T����N��N�cB;��*����wOx�Ny�ǥc �auu�t�ERM�$�&���Y   � �a#ɏ$�V:�"q��R�.�W�n����'��F�Yٽ�����tD ����#,��$ߗ��%y�p  `�)�  �U�|W�O)d�8I�y��j�B{��I��(	X`�j5����>�A��nvvv��v3' �
y"�'��I���   L�  (��%���!��� ��J��V�����t:�,//��gj��g���$�u:��j��0��z��׳����x����Y�}��+ p�g(�&yg�/-  X\
�  @I_��ϗ�����JG �9:�}ee%��C���x4�pg���8�����3�vg�L�g4���������~F������f��[7��I��#a�lo�?f��=��lo�3�Y�^O��~�}�'\�X?���I��VVR�V���tR=,��z_����v{V�-/��lN�7��^�R���|�J���u�\k�S��OL/�i�Z�~�z���쾳�c�; �#����I��$__:  ��.��c  `Q|f���R:ȢRp�q5�ͬ��dee%�v;��_�gaZ���L
�;;���{{�z����������x8����ϊ���-�O�ݣ�݌����2:8(���x0�`k��=q��;�DgoV��TR_YI2)ԧZMmy9�F�X�q���n'�ZjKK�.-M�?,��:�T��Z�T��&?��J�јl�VO��$�Z-kkkY[[�x<�����ׅ ��2����M�KI��t  `�(�  %�)�$Y.d����ÚN6^YY���j�����`{;����`k+���;��~���w
��nF�A�;;�"s�7{���x8�`kk6u|t�$s�lF��)�o���V'����;e����Z�T��YѾ��6+�ז�S]ZJke%K�zvG�����'���r}�ٜL�w� <�V��F���]w���T��#�/gRt  87
�  �yk&��$�+dљ�����j�t:Y]]���J��j�H�dtp�a��a����V��ެ|>�ޞ�lOZ���po/Ý���&��#�v`��F�I��[�%�=|��N��aٽ�nO��G
����Ia�p�}��J��Jm���N��N��u�p X$����y�f��l-�{�|z�!  �s��  ��o�������� �5-�O'��,��4������v�������ome��u|����d����J5I��1Τ��K���g��g����:�_m6Si4R�t&����T��f��k�v�N*'�wX��	� \p���
��}r��M�I���   B�  8O_��+K� �V�i�ۥc p��j����dmm-�N'��(=�4-}����wv2��ɠ�ͨכl�ٙ���s�0o*I�Ӳ�t��i4�F�~F�����Tj��d�Ng2M�՚=���;������]Z��M����������%��$�t  `1(�  ��O&�_J�`bmm�� \�z=���Y[[K�՚�n�zw��oo�ylme��3������t�ay}���a���`P��\G��9�����t��=]�R�Φ�W'�O���_��k�S;�0_�tN�� pY������1�J�/
�   ��;  p>5�?OR-������ 8c�~2�p���ͨ��xw7��0����z������E���n�Ψ�/�ҹ��~����Qv��hrW���Gz�ѸS~��_?,�O��G��WWS�;�p�9�u�T���$L�g  .9G�  ���I�t8� ������e��;+�����^F��d�����p�����po�؟UM�J�N����*� ��J&/��d�i�}T0W	�~?����77���VkR~o�'e�Ng��#    IDAT��p�zd�|�p����� s�1����=I>=��   ���;  p�*I�'�o+������L'�vv2<|�,�6{�v3>�<�j&��i��r
���wt��8��{7����`�y0���pw���W�VS;,��WWg����kw���Zg�	 x-&�_HoH�%��$n�  �	w  �,��$_\:�rr��L���^/���nݚMP��ܙ�~8i}���v2>���R&�OieRr`~-��2)����ڛxh��(������}�N'���cS�k�Τ ����]�I�%f �Ð��3���$�M�   ���  ��/I�5�Cp2�w�Ѣ���>������[���[[�F�����I����V8 ������$��)��������J��+W���H��Q�x�a]h.�/%�{��   ���;  p>%�w����w�2�log�����v��Y������_��dԟ����3)�w� �eWK�r��'�fRv��y�R|��L}uu2~m-���IA~u5���ɺ����j*���%g����MI>��J  .�  ���I�$��p
��Evt�zs3�[�f��;;�u���������NV?m�$˙�[��X,�L�����4�n&���%CqjF9x�����_m4�8�_�t�,����_��Z�u��N����<��tT3��'��$�^8  p�(�  ���I~[��:�w�Ӹ�Os3�â��p��tݰ��p����wwKG�p�\A։ۣ 01��i9�I�Iv2������ٿq#�7n���F�%�z�����������h��j��땎��]O�/���${��   ���;  p��!ɗ��ks{g�Q�����3���`k+�۷3��N�����������GS�dR{'��; �O-���� ���$�qԨ��hs3����ܷ�h������z�kki��M�76R��Hcc#���4�^Mui���lmmM�����I�E��,�  �$� ����I�f�<܁�����������͌��ܺ�a��a�wg��V�#u��2���N�:| �y��Ȥ�ދQ�<�Q���͛�߼����=~6���<\6xTkkky�J�ൽ-�H�-��   �O�  8�����o��0��3py����LW���`{;��������o�����x8,y��2�Ծr� �����N�A&SݻI���=�d�j�1��ʝ絵4�^�L��r%�É���Qkkk�#��)�/$���A  ���|  <�f�Hr�t���0߆������ܺ���f�_z)���72�vK��-eRj7���TO��d-�n&EwS�9o�~?�/����_~�}��l�ѩ�Ǟ�\I��T',ǲ�J=�w%��I��  ��>  ����$�^:�IA����q���߼��[�ҿys�����+�L�o�ʨ�/��TM�Τ��(���R��wP;���;���G%C�	�n�n��{�U���������k��{���I	���4�^M��`�9�5w^��@�?7�  ��;  �8�l���t���j��pƃA��ln��p����w����R^y%��Y3�R{;��P^=�F�Lu�N�2:��`k+����~���ݧ�h���ө��+W�|��;��]K�Z=����Pp�K����&�K��   �I�  xToN�J��᭯��� �ʸ�OssVV�>�߸1�Ⱦ����_NFf�.�j�V&��f�, p�j���� �����1����F�o�x�������a!~�p]���TM��"k�[!�L�]��   �G�  xk��f�S:��+xp�^/��7'�[���f7o��֭��J�ne�햎�T���j&�A ����z&E��$��������y�U��w:�_���իi\���k����ki\���k�./�SbX�5̭J����M򋅳   sF�  xX�$�N�J�јz�nw2q��i��	�/��A�W:&s��ɴ�v&�0`U3�Hk%�n&E�����bt�t������O�ј�ߟxb6���w&�_�����9���gX�\�$��$�'���   ��;  �>����Spg��ܼ���/g�p���+����sp�f�ne40���Qɤо�I� .���v&��${I�%C�7����F�o�8y�J%���;S߯^M����T�k�Ҹz5�����rI�r,k�}j��H�奃   �C�  x(�ה��qR�y7���OZ�q#�/�d�:箖�(���e �̖�LƯv��&�95��$���]��zj++�I����+W����.âX]]M�Z�h4*�G�eI��$�R:  0� ��d�w&i���YYY)�k<ep�V�_~9��i���7s��+��J^y%��;ZSV#�R{'�ɶ �H�I֓�%�e2ս_4\>�� ��|�gNܧ�j�y�z��x"���'S�_����_�����9���S�T�j��u<`��I~.�ϗ  \|
�  ���&��$o(��g�;%��ɤ������b^z)/����l\P�$��L��EW��b�N��L���E�b��f��g���'n�6w&�?�T�old��'���i^��T\���X]]Up��$ߛ�w&�U8  p�)�  ��|v���9K�~?����߸��728�:8-���r��Μie2��Y: \P���A��$�Pިߟ��l���g{�^O���c���a�}��'Ӹv-�j�@r8���j^x��1x|��I����g  .0w  �|Q���tNG�ZM��)�96�2x��%�χ���ۥ#©�$igRlw  L3��L~�>4��b��I*�ZW��y�z��xb�|X�o^��ƕ+眘E玄���'��$o/  ����  ^͛�|{#�.�N���[����~�ľ��s��g����d5I�p �W�$��>��d��{��|���_z);����l�N�o>�D��zjR�����SO��nH�e掄��7$��$��p  ��Rp  �{�\/��c�S�^/�/����<{�?��>��)�]-w�����Qˤ辖;E�a�D�i9:~���g{�әL{�����i���<Ǵ.�z�w&�]I^,�  ��9   ��[�|V��.Ӯ�x<)<���������ǳ��g��U:\�LJ�$�o g��d=��{7����h"����y&�g��g[�ZMcccRz��4�z*KO=��'�L�u�K��*����1�K�u�X�ܸ�  pw  �$_��ϗ��s2�r�����ǲ���MJ��?���</���@uN�Ȥd�. H%�J&���lE��x4��͛9�y3;��+�l���f���f���%��)���K�s���$_[:  p�(�  w��$ߞɐ=.'�_�֭���},�g��,?��";< �v (��IɽEw�^����lo'O?}϶j���Of��o����/=�dׯ�Rq_���1�K�'��$��t  ��Pp  ��&��$WJ�l88?��������{���~�����_Ϡ�-�R#�j&e: �b�ݏNt�M\t�~?{�=��瞻g[�ٜL|?�������
��������֥VK�Iޜ���Y  �B�  8��$���!8;+++�#p���t?��t���}����y&��z<.�v �����0�F�}���>��=۪�z�O<1)�?�T�^��,=�T�_�z��9�֥�d&�W>7ɸp  �Pp  ��0�_*��e���q��K���f�C�ί�j�>��d����F��L�r ��Pt��h0����g�����V��Ҽv-�'���ߘ�7�i2����1����$_���s   ��;  �$�O�I���p��<?�~?�8��>���O���2:8�pw7/��A�W:"\J�� p9(��e<f�ƍ�߸��~�ضz�=�����O��o|cZozSO<������t:�V��F��p��!�O'���9  ��� �J����6�\rn�|�F{{���Cn��ϥ�k��Q_�K#�z�V�  ���ݻ��e� f��e𑏤���[_m6��������4L|?3�J%+++���*��UO�]Iޜd�p  � w  ��|^����Fs37~����O�d������B����v5 ��:�3��v�a�8�����3�=�̱����,��i��MY:Z|�v�P��E�}a|B&Y��t  �w  Xl���o���1��t�����������/����q`�Ԓ�&Y�b; ,�J��w2��>*����^z�HzwM|��Z�I��G�W�J:�nX(,�_H�J  �Pp ��u5ɻ�4J�|T��t:��1.��G>�_��o���ϗ���I�}�p X<�L�t�lgRvWt.���nv�~:;O?}l}���շ�%o�3�P����p��$?���)  8� ����$o,����tR��s|n������߮�稚d-�듬�A- `�}`=���.�|t����_(cn(�/��$ߝ��[  �c�;  ,����J��|9	x
��<��w�Ə�X�$�0*�Lg]KR+� ��jI�d�}a+I7ɸh"����K��l��r�9���~s���*  8_�] ����I�^:�oee�t��6��w�C��Q;���W�� ��i���$˅� <��h���+c.8����*�Y:  p�Lp ���L�L��`�|t�?��|�]���/��a)���3 ��j$y"�^��$��q ^��sϥ�ɟ\:ƅ���B��$�O�L�   ��Pp �������t�p�7���3������_.B=�Z\� ���L��Mr;ɰl������r�t�9���B[K��I>+~� �B��   ��?��-�r�|8��<�_���Sn�sP��L��� ��N��'وc�Ŵ�쳥#���g$���!  ���8  ,��I�Y�`�9	����>O�7�����Q�R�$Yɤp�~� �,T��frA�J|� .���+a.�@��I�9�C   gO�  û39��s��wv�o��z��Q�R[N�T�+q�
 8?�L�<��������͌vwKǸ��"�_�ߙ�u�  �%��!  \~5��AyN>�����ٿq�t����ʞH�(� X\�L��\��$�0g�c+���k�Z���cP�'$yG�  ��Rp ���w'�[�Cp1�����p��~��y���/.���R�
g �j�]e��a��JG��*�J:�N�\_��K�   Ύcu  py-%yW�u�C&�����ތG��1���$y]��$��Y  �V��{��2��P	���-���$��t  �l(� ���-I>�t.�_�pw7�?���1�RYʤ(v5B _-��-O�g����@�9b%�wg�+  �d�[��g�΃$�����'�y��*+��2�>zfZ3�:G:-����&8���#K^H\���]�»f9�?�`�]9 ��� )4BB��cFs�Y��u��GfUWOWwWwg���|ޯ����|���ROW���<� `8}�����p]�-��b�ӟV�Z����rXQ�g�  �^�j�3.s ��	��C�/򤤟�   ��(�   �g\��qJ:���8�1Bm��_�� <G҈�S۹�  ���?׌��s �RmwW��=����8�?��F�    ���   0|�����[���3�XG ZBҤ��8�  �����7EI�q ï|�u������JJY   �=�7   ���$�w�!>L���V���ښu` �%MH*H�   �v�}\R�8��ut��u���n�I��:   ���   �I��u��wVY[�Z-��@q$�H���4�  �/i��a~0�^�0������;�!1�   q�     ����F�� �X����Ɔu`����:� p,�L��n���d�8�$ɉ�K�O^s�@���|�۞�⸮�.�s|_n�|O����>?9�LJ���%7���=V�ۻ��t��=��rLc���N�VS�\�$5�u5�/4����wj�x,�^*���8~��/5�w�+WRNRJҶ��m C�	�w�9.܁#�_I�I��   w   `8�G�߰��b����J\ n�U�J��ګ� ��tQ<���K����r;E��8��DB����}�	�q���r�qqۉ����S_�X������hk�U���<n��jV���f�r�q�z�h_��qt���N��V*I����j6jH���j��j�|�f���ڧ��_RQҁ�]I\��A�)���pE��|�u    ��;   0�^!�}�!n�SSPq����R ��R{R��g&�K��z^�>�A�X�+�J�L6������TJ�����N��ssy=����@��R����l�0I�`�)ͷ�uՏ�����4�ە���'���}��@�rY�rY��=����#)#)��4��m �����Ύ�\�:Jhq���~Hҿ�   ��Qp   ���D��:�VwV/��# ��4�viT�﷋��t�P�%�����y&Ӟ|����=�}|�T�fO��N1=��7��0 Lbɤ�L��h�j6���o��e5U��o?>U�ot
�����㣣%�r��9GG�׸�r��%�.�oK���0��׮Qp��q�>$��%=o   ����   �_��r�?��l�_�� ���4���c��b�����X:���ȍ�y2��Ȉ��t�q���dڟ�J���dK����{ @w9��x6��"�M��K��Ǎ���t�NI�V*����W�s�88P}�}�L�G�%$MJ*Iڗ�� �U���<�u��J$�<O�Z�:
�-#�$�E|;   w   `p�N�OY��``��۫�J:|�aN�i��S�=� 8��*�ɴ���l������d�v���L�]<�|K���u���� @��i�����������|�vR���;y��������;�����Zu��WRNRJҖ$*� �Eyy�:B荌�hkk�:��Mj�?��u    ���;   0��'��=Ĺ0���v?�9��M�@(���j�9cj{4�TP?u;�s�i� �p8���/��k4+��S��OO�otn��]���T��U�s߬T��'<�����%�� Χ��b!�2�w��/I����b   ����   �_���Lp����>g�@Ҹ8Y4b���\�d��I��%u
� ��� �R>_�߬VU?�����z~X.Bu$�HJHږ��?���~wr�=HJ�CI���0�   ��f	   �7I���!08\�U���Zͦ������:��N= |�x\��⣣'�Ǐ�\��s�l���y�zl� ���
��{����ލ�{��Z����[�TR��GG=��<8ORAҁ��܇������j��r	�(�E���5��#���    8?
�   �`II�=�<�A:���8�1B���gC[��������~{���T�ν_(ȟ����*62"��1^>/�u�� `�xw�`f�?�^*���q�����Ɔ*���"����}u}]����	n�H���4�r_���i�TY]Urq�:IhQp�}�YI�����   �|X�   ˇ%=b��E����җ�# &\I9I��p�XL��X�6>.|��8�k��s�vI���u'�� @d_Tv^��#�wwU��Vu{��xg�侶�ݾ�����Z����Ӎi�;b�;�[���)���p|I �U�j�Y    �w   `p�7�~�:O&���Z{�A	���S������(����������r
&&?.���+>:j  tQ,�T,�T05u�ϩ�﫶�uS齶���Ύ��B|}gG��Mն���9*���:Ls�b��e��ƹ.ܧ'$�_�{��    �;
�   �`��o�����֪�t��3�1���IUt����2�՟��?1�x6��P�?1��Ȉ�lV~��`rRN��d  ��♌♌��<�Y������ޞ�����V*������ummmimu�=A�TR��\w �*++�B�s]x ?-�O$}�:   �;c�   �4g��m�϶����YcGbDCRҘ�1���Mߤ������(   '\ߗ_( qF    IDAT�/�z�3��V�Z^^����j���Ƿ�ݓǵӏwvT����`Qp�3�u��%����K�(   b�  ���FI�o��E��~�k���s՞���v���~��)� ��������]W���>�Y.��ݏK���v1~{�=5~kK�R�2<0 ����B�s]x@�Iz���X   p{�  �p�H����(��m��v@�C.�4�h����S?%/���  �@��ǕN�u��u����&
��LM������j;;����ꥒ�����v������Gp�GG����B�����.�'��/I��   �lQZ�   �oJZ���Ƣ��(�cX9�F$e;��b�e/S�[��:  @WA���%mllhssS�V�+_7�N+�N+1;{��Z�Z������ޞj�%���wvT��QugG�RI�z�+� ܬ��L��68ׅ.�$���WHb{    �(�   ��vI��u>�nU]_W�T��t����v�:�����.ɉR�  ;�qT(��dt��uU������������w=������n������������R�Ύ�������h�!90<����c�Y�%���*��u��%�O��Z   p+
�   @8%$��$�:_&���:�<c躌���5��X�u�S����  ��dR.\���vvv���">2��Ȉssw<�qp�Zg�{}{�=��~}�dJ|���Sr �*kk�Bmdd��;��g$�����   �f�  �p�����C`80��V�>k蚸�S�� �~臬#   ��뺚����Ȉ���U�׭#ݳX:�X:����m�i�j'%�Zg
|mkK��]U77U��7�8��R^Y��j###��ذ����K�=I���V#   @�Pp   ��m���u&����k_�� tEJҘ���G��4��W[�   �L&�.hyyY����q���<����B��5������4��榪[[�u׶�T��}-U
�w�@t��%�O�~�:   �(�   ᒐ���vW]亮��u�Pi�j:�|�:�@\���)� !0��wZG   �x<���y���jeeE�f�:R�ŒI�fg�7~{[��U��T=~���~~wWj���8���Z���XG	%:���+�����     �(�   �����J��z��^P�^���7�u5��+5=���v��T�޶�e"�J��-�b  ���訒ɤ�^��J�b't�3�U��L�om�ڹն�T��Tu{[���>�nh�˪����嬣�wt�/����:Iѻr   !
�   @x<)�ǬC`���w��g��� ܞ���?>.o|\~>//��76&?����k��G��o����7~�a`[�o~�b)�� ���}_KKKZ__��֖u���x���)SS�=������*��nn����~~cC�j���%��
��9/��k$���>h    w    ,\I��Y�pI���B��k_�����ӊ�r�r9���r9�s9Ţ�\N�Ą� ���b��fffnY�///���ۯ����ۭ#   �s]W���J�RZ^^V�Ѱ�4T�S�o�����Ύ*kk��������Ύ���nl��d 0�]umMz�1����bg���K�cI/��    @�   ��Jz�u
�:|�y�R�TJ��q���	��S��ޯcJ�Ӛ��Q<~�i�����F�������&�   �122�D"��ׯ����:N���i��i%fg5����~2~kK��MU66T�ظ1	~cC�Z� 9®��j!����IK�7���   0F�   �����X��pb��f�rY��u�@���/䏏��?1!?��76�.���r�����8���*
�=��_��{��K_��   n�y��������8�8��z��.������~r_��Pu}�|D�WV�#���Co��j�   ��   ���$z�	�nV�rEj��c �\�k���

�Ţ�\��.��[��433s�-����>%
��+^a   ��Q�PP:�ֵk�T�׭#��٬�٬�.��z��@յ�v�}mM��m�vv�e���ըT���Pe��m�k!z�7$�GI\e   ��   ��Q��)z�����\�� #�+����{Xd�YMOO�uݻ�	��  �(�J顇ҵk�tpp`(�N+y�¹��uUVWOJ��j�ω�������}��zPp�=6&�%��    @TQp   �LI�%�nw��5e
�C+�N����-vrR��o�x�f>�?�����v�!�R/ZG   �X,���mnnj}}]-v�Z�[��������V����8�F��Z�$ot�:J�PpG�m��l   �"
�   ���MҸu7�nvt��u�'otTA� obB~>/ob�]^��;�o�x�����{�(���g{�(�\�Wbr�:  �����J&��v����u�S��h�������j������I����ݞ"��
�gH��r]WM.�@o}XҟI*Y   ���;   `��Hz�u�t:m!Tʗ/[G�m��מ�^,�/�����bQ��YG�t:���Y�b�{���K�z�(�33��Z�   (�TJ.\еk�txxh!��b�����j5U77O
��UU�������(���8Z*���<��u��qG�dR�Q0ܦ%����   Dw   ��2�>d�@����֖�8Lycc���z�s�
�r9�x&������}}�ѕ+]N3833�   R<����׵��i��<SS
���|�V*��)����T��kk����9�𩮮ZG�t:M����%�����:   %�  ���uIs�!�L�:Bh1���\߿i�_,*��8yn���߫X,�����%��c��  p��Q�XT2������u$8/����*}��-�5+����WN�߫j5��Kye�:Bhe2���Y���s%����I�g   "��;   �_OJ�!��
�7Dy�u7ųY��JLM�/N��^�(ot�:�@H&�����������V�7���   0�FFF��^��J�bC�%�畜���V�����M��ӏ�����;���%����X   ���;   �?Ǔ^�9}�8�M�6����f�wJ��Ԕ�bQ��I�SS�%���Z.���Ԕ�y�U��6�T�:  �P�}_KKKZ]]��ΎuD������5r��������U�~����'��1*�o��;�콒����Y   ��b   �?�T�+�C :��\׵��o�e�
:�`r��LMɥ��u�XLSSS�f�]�����m  ��u5==�d2���U5�M�H�$��7:��ŋ
ff"[po�˪��k��>K�=����A   �(��   �Ǽ�n���Z��*���1L���Mʾ�U���$%�>�}_sss
���_7�����u  �����H$t��U�j5�8�M��I���������/x�����9   ��Ǹ+   �?~G:s�e�g�buCyyY�F�:���7��^�z%��(��Q:�օ�^n��V�'kRp  �D"�.��$B'�N+ῗ��U���J��# �>$i�:   0�(�   ��NI�:��B��+W�#�r\W�������5??/����X"ѓ�;�  z&�i~~^�|�:
p?�S�+++�Bid�y"01!��!   �aG�   譌�߲�hb���ׯ[G0�OL���q��u]��̨X,�q������=��a�w  ��rG�bQ���=�`�WA��Lp?�`��Iz�u   `�qF
   �!i�:��E���t��㟡~�}_KKK��{E�����u  �H�f�ZXXP<��D�����ù/r%�+I|�   z��;   �;����C ���~Cey�:��$��H�RZZZRЧ�y,���ʊZ��u  �HH&��p႒ɤuD\P,ZG0���q����3�!   �aE�   ��\`�)Vm�V+��Lp�\.����b���g�'��&  �Q<���r��uDX05e�L�\V�T��:��4o   F�  ���QI���hc������f�j�Tbv�:��rG333�����8}}�(�%����   ��8����M~�$)����`*��%�N����%�/�!   �aD�   �1I�0��-�S��Ubz�:�P:�b9::j��n*e�aqt��u  �H�ؽ��x6�X"a�L��o��u]%�I��wH�N�   ����   t�oH*X� (��U���#�
���x�u������L҃�	���2w   3�TJKKK
"����/�#�a�����!�[���   tw   �������! ��c�O8K��ZG:�tZKKK�/��y���V�r�:  @������%.�F_SS��Pp?���~�:   0L(�   ��H�]I�эP�d��-�ss��J.�����\����7>n����O[G   �<�u5??���1�(����u3����/��OKz�:   0,�Wc  ���^i8�����uSLp��q455���i9�cG��OLXG0UYYQ�T��  y�?+OF�x��	"�����f!�8��	$}�:   0,(�   �Q��s�!�c����<��Z������1L%ff�#�X,�����M��y�����U�   �����b16�C��Ţu3��5�c�w���%}�u   `Pp   ��7%����Hcq����*5��1�8���ۻ��}---��)����~�:   N�d2ZXXP<���!LMYG0��[��i���}HR�:   0�(�   ��u�0�q-����#�������u���J����$?�����1�   |��.\��D"aC�����w�~���[G
��YI�   :
�   ��q$}X�l��aq����b�T0=ma`���jaaA�X�:�m�A���uSLp  �x<���E���XG��q�Ţu
3Lp�CR�H�c�!   �AF	   x0?&�5�!�cq������W>���̌Ǳ�rWɹ9���^�j�:   �ຮ����筣`�$&'�#��Pp�CR��i   d�  �����s�!�����v��l�T�	���qMMM�8@� ����L�����1   p�bQ�.$����}���[G�< ľY�wZ�    w   ���I��Y(��U">�����O���rO/�KR�_��   �����\��I<8�.J�*�oA�!�[��   � �,   p�����C �C�]j���g�T05ea �b1����x�'�K���h   ��f5??�X,f.ʿ�V66�j6�c�
��r��~�:   0�(�   ����[� ng�����f�����c����ZZZR*���r_�ss���~�s�   pN�TJ����<�:
X"��[��j���1B��;��%q   �G�  �{����j��d2i�\u}�:���ԔǱ�j�dRKKK����^)���֖�ׯ[�   �9A���%%	�(P�Ą�x�:��J��w�X,S�1�;IK��u   `�Pp   �MZүZ� ��UR%�܃�i���N�����X,f���㊳c�J_��u   ܃x<���E~w��q���u
3Q߱�,�[��%}�u   `�Pp   ���K���M��k�'�SS�B+��i~~^�;�E���Qp  <��j~~^�l�:
P09i�L�w�;w G҇%��   ���c%   菇$��u�<�ɤus��/�&��~���	MOO�q�(]�~����(�  $�q4;;�|>o&����Xw
�OH�1�   ����   �߇$%�C ��������399��nc������V}o�:   �S�XT�X����G��^������R)��y����u   `Pp   ��풾�:p^Q_�k�Z�nnZ�0�OMYG�q4==���q�(=�wIͦJ���u
   <�|>�)~��9%"\p���g�d2������   � ��   ܝ#郝{ ���b��uS��5k5�f�lV�d�:F(8����Y�r�;+}�u�P���g�#   ����ivvV��)ܙ����}5���c�J�=`����ǬC    aG�   ����j��y��'UVW�#�
"<��4�u5??����(=卍���c���  0�٬����,c����	9�;R]_��*�t�:p/<I�   �]t�   �'-�}�!�{���,�Fy�ݱX,�����,r3�]���W�88��  �.�d2������d�='W|�w꺛�_��bQ��C�[$�M�   @�Qp   ������C ��	�R%���Op���Z\\T2����7ܥV����?o   ]�J�����x<n!
��T�֬#�
��0�>$�or   �mPp   noQ�?��+�X�MDx����Z\\T�Q�*��#�Ba�3���   �.
�@����}�:
B(���Q���Ř��uQҏY�    �;   p{�%):�142��usՈ/��]�r�%����Ba��;  �Љ�E��;/��#~���(�c�����u    �(�   g{��wX� �ܥJ�'�SS��.�JiiiI�x4wvN.-)Ƃ����%����c   �����H$�� D��	�f(�ߌ�;ظ�_�   �Q4W}  �;s$�f�8Q/��j5�vw�c��%����X��t:���9�nt��w\W�G��g?k�V����|F����:	�ЬV�,��8<T��P�VS��H��(�ժ�ڏ���j6�j6U�ߗ$��U5+IR��P�z�}l��V�����-��8u왙�e5;�{�׫�[���Rr���X2y��n<.�E?���i����ǎ���L5�%�r=O���M$��b'@�29��~�sL,��G��@�� @�b1-..����:�|_@��Q�ྱ!�Z���K��;�K������    aB�   ��Hz�u�~e:������y#*(�#���F�x��������X�ZU��@��C�K%5��ԬT�88h�v\N��T��W�V;)�7�u�K%�����u������s�<H���ˉ�o��;���i�(�����(�H�M$�d�&��ǩ�b�̍�FF��DB��_�	�������]�zU|ψ����{Z�VSmgG�ؘu�P���<_�Ŏ�   �M(�   7$��u�AD}Q/��t������r��F�x�:B(�|�S��Ъ�����q9��@�����>nt�;>��y���;M:�ph��j�˒��ϭ0�T�]v��>�&�%�e2�w^s��vi��Z|dD�tZ�ų���##r=�G)��뺚����������jF�g����������g����6I��   �w   �f�TҢu�AD��^Y[��`*��{&����,��S2/}�u�P8�tI��U�o�ӬTT/���RI�RI�����O�~r���t�J�s1E7
���+����ApR�?���Y�FFn�?~��g�4��!I�����U^]��b�����ŋ�1B#�NSpǠ�MI��ݭ)  �S8k   ܐ����!���d�#����B�:B�e2����q�(�����76����us۟��������f����j;;�mo��;���wvn*�����c�ԬVU�ظ�Ϗg27M����3�s9�cc�����˝�;\h�r]W���v���Y~�݂{���X*��6�c��J��H�#�    @Pp   n�%I��!��	�/�OMYG�l6�����y�K���[�0���S��_��-%�����Ǐwwo<��8:�N��������=����Tx����W��7:z��W,��Az �����,%���E޷S{����Q���"�%U��    �(�   m%��u�"_p�ܴ�`*Q,ZG���QMOOSn����^F�]��SOI����<�V������[[�nl����������������mȋF    IDATm���-5�֑���-����7⽱1���������	y������
�%�=L������U*���ςܙ�~���h��1/�]�~�:   `��;   ���|�@7D}A/�w��������'��WXG��֖��yF����:
B����.�������.�oo����PukK��U����2�z����9'�ƒɓһ��˛������

����z^����8��NO����q�G^��Lp�Y�>`��G��J��IN   @�   I����:���ɋp��U���m��Ba(�\N����1���}��x\�z�:���O~��{��vvT��T�S\������yRd?��Y�YG�si���]�r�c㣣���v�PhO������+>6��Xl���bH@j�܏o��Q��^��T���� �#�N[G �%+���~�:   `��;    }P+A
Q�VU�ܔZ-�f��I�]w<��K&�y�Q����j����?�����f���ꪪ�몬���'���4�f�j ��wwU����s���8���ML((������bQ~�(b���XǓ�%J�Q�G��ެ�T�ّ76f%(�c����ߒ��u   �
w   D��Hz�:�-Q_̫F|{�X���U���'��_�����.��/����x&cwЬVU]_o�66T�vM�S����mm��lZG��ЬVU�~]����x\<�mO�?�
J��ʟ�PP(�<�����Z��J��u�X|dD�DB�r�:�������}���$����e   �B�   Q���!�n�|�}s�:�)�
��l����)��W����us�z];O=��o��(�լ�T]]UyeE����_WumM��$������  �ꥒ��'�ǒISS�{��`jJ��)�[bfFn�15p��I�܇�_(����&���J_�h#�~NC���,�/��    (�   �~\�#�!�n�����֖uS�2EsddD333r�:�@}ի$ǑZ-�(�?�I
�=ԬTN&�]�z2q�������u Z��#>�����ǜ����Sbv�d�_((����}L�(9.��Z-���Y�AQ.�G|'��(�c9�~]���    (�   �R���u�ۢ��W����	�lddD��������)����^��bn����0�껻:�vM�k�T�~�=��3��������uD @ȝ����S����337��OM)��>�8(��Y���sG����z�������G��b��Q]_��Q?'������]��c   �7�
   ��-i�:�mQ_̋��`����4��.ɾ��%UVWu��J=��u�PjV�����:�zU���U>��N	 �c�J��S�]WA���쬒�����̍I��|c 9����9J�C,��
�Q?'���k�>*�-�   )�  EyI��:��T�:��(Op�g2r	��-�Nknn�r{�����Z����:F(l}��.��K%�;S؏oGW��//KM�� !�l�����ʊv?�[^v}_~��.��͝���J.,(F��'���Љr����O��91��%}���3�   �w   D��%�Z� z!�ӪZ-U���S����r���Q���OZG��O|Bs��}�1z�qp�.�w��/��ެV�# �3�j��������u|������Y��J-,�/Ò뺚��ӕ+Wtxxh]4ȿ?���Z��K�d2��^���'�b   �
�   ��I�:�+Q.��J%5k5�fuA?�JQnXTrqQG�.YG1W����8<TlP���Z������e]�rRb?.��ww� Zխ��E�_��-��A�����J��+ٹ%��P~Z��j~~^�/_��ёutI0��wC�^W}gG�ؘus����<�"|nCmN�?��A�    @�Pp  @�����u�W�ɤu3Qߖ{��ɤ���)��H��.�Y�i���J�o}�u�;��J'h�{N�=�.�_��F �f���g���3������%fg�z�!�zHɹ��4��i9��:�\���.]��r�l]�&�g2���[G1Q]_��ޑJ���E�^��I%�    @?Pp  @�|����:�KQގ���e����[G�'APn��k_��?�c����񏇢�^��R��^���ի:�|YG�/�|�*%v  B�Y��\x���S7�K&oL|_\TjiIɥ%����Z��tɽR�X�A��b��闼�:F(��i
�f����w[   ���;   ���$ŬC ���p���	�Ţu�s�}_���'��rO>)�u�j6�����˿��{���~|;x�Y>�ld7  ��ё�~ZO?}�k�lV��~�a%fgO&�'����B�XL���t�j��u< bB��=g�De}�:BhD��"��%���U�    @�Qp  @T�I�7[� z-�LZG0S��wb�:¹��q���+�D��GG�~��Q������^��������.]��K::�]���+WT/�S8  QU/�T���U���oz������pAɅ�.\�Fi!I��Lr����q� ��n�Rp?A����~I?b   �5V�  �"ɱ�Z&���`&�����Ŵ�� ����D��ORp����'��^/�t��s:xi��=��^���  ΩY��v�?1��C���=����*዗��x��K�.��hX��}��f����B��;"��ޭ�Y�    @/Qp  @|���X� z�u]%	�f����fC?��u]���)y�a�{�ku���[�����k�{�����)�.���N���I @�T76T����SO�x�u���U�ᇕ�p����r�X�'� ����._��&2� �w&��H�R��~�$����   �w   D�/Z �!�L�q��QA��a_�wGsss,4}�k�z����us���k�|�S:�z�]f�����++jQb  a�l���]��͏}����ܜ�/�o�<��ŋJ��H�]�[�ɤ���t���Z-�8�G����j���H���~Yҗ��    �B�   �^g�(��[���{{�1̄y!�q��̰�l$�Ji��/��g>c�\�Z��ǭc   ܿfSG�/���em����<K��\\T��e\�V��Eycc�aS:���̌�]�f�����n$/^m5�mo���b.���9�ڃ}�i   �
�   f�����K���ie�OLXG����)e�Y��6��7Pp  b��C�������я�<���Q��G�y�1�{L�����&�lV�FC+++�Qp�S<�Smk�:����&w1���^-��A   �^��  �a�}�^n�H�77�#�
�E�g���T.���ycox�^��߶�  �>+_�������O���9�PP�Sv�<��2�?��',�����hh}}�:
�AP(D�ྱ��ŋ�1�%�I�@?��~E�7[   z��;   �U\���C ��E�Z��a�����5���Pȼ�%�'&�;    Ҫ���Z_��_���s�Ą2�?���W���T��/��H����	5mE�0=���	�_��a"��E�Ey�"뿕�fIi   �6
�   V?,�a�@?Ey�J�a+��������p�^�:�}���I   BՍm��_��ޝx\#O<��7�Qcox�ҏ=&�u�Sژ��T�����u�C09i�L�w�;F��+��b   �6
�   F���X� �-���Q.�;N�
��tZ����1�"c_���  p.�z]��^��^/������{��5��7j��oV|t�:b_MOO�^�����:
�"L���6
7�=��Ϭ�    �D�   ��'$�[� �-ʋx�ܽ\N��Yǐ$%	����q�(x����z9��V�i   �����?�S�����<���*~۷i�-o�����z�q����^P�R���;��f(��E��"�E�   C&��	  `�����u�B������!�P�y����亜j#o|\����  �׬մ�������w�S��-z��Veu�:VϹ����y!��g�E�fj�B!ʻ"�^#�ۭC    �Ī3   ��OJ��X��"^�'������({��[�j   C�^*�����>��w�+�}����%�H=��5??�X,f�ፍɍGs���GG�1���q��Y��_�Ķ�   �  0LI�XI���L4+��c����jnn��0���XG   �j5Z��?��~�����i>��u��	�@sssr����8�#[�2�]R�w8D�}��wX�    ���;   ��?��aQ��^�޶�`�z����4��"}񢂩)�   V��6?�1}���[_}��T�~�:QO�R)��p�)���	�fj���B�s���)�   �  0,��@dEu����p�~rrR�l���q�G�o~�u
   �V����~T�]ߥ����ժu���f�*��1p� ��#~~�XTϏ_'�oY�    ���;   ��O��툸�.�ՙ�n��|^���&����[�#    "���.}�#��w�v>�)�8]��D��	�[[�B!��ǀS�/��  `Pp  �0HJz�u�ZT�/������Q���'�T,���  �9�|Y_����������q�jrrR###�1p��E�aP�ذ�
Q=?��2I�   <��u    ��%i�:`-��j�'��	�2���g"����T_�����r��6?�1�(x@�Ȉ⩔�x�����J��x\����f���ё$�~t�f�&I���~x�f�n�  DR��������O��_�Ee_�r�D]333�˗/��sl�Q.�onZG
�$�$����u   �~Qp  ��KI�I��5���y�u���=���<����u�n����V
�!�}�gg���VffF��I����y�cw}��Ͻ��j-�$�j��mc��`�mC�6�� `[� �2�0�$3����0���p29�$�2L�	�<,�L���q ����^��k_�>Twu�{�E�W���:G�dI%}�������/Q((����W��)��)��/�	+KKZ������ssZ����쬖''�t옖��ұcZ��k  @Z=vL��ַj��߬]oyKS��X�}_��㚘�P��	��XG0S��.�����,�U�>g   �.
�   �v����荒��̴s2],Ӯ]�J�v�;���j���Q��yʌ�������u�^s�F�=��2N�N+L��7>~��U���x�����¡C�}�1�>���T�\nSZ  �+��}�SZx�a��)h�T�����u��!�y�m**���S��V�^�Gv�	���#�/�w   t)V�  ����c�./ޭMMYG0�΂�����x�^�
��t�~�:J��b1�o�AśoV��땻�:�_w��.���R�_���_���Z�\���G5��i��I��E��  ��L�z�o�͟����w[�ٱD"���Q9r�:�Ӽ0T�ͪ�����z]ՙ�����i\<�Mb�;   �w   t�wI�tW�jU5���a�Ж�R��*��]wQpo� ���Ӟ�ҭ��p�*=�z���)�o�r��i�K^�q��ѣ:����C��Ci��A���8  p��Ç�Лޤ�~�w�{ֳ���X__�599i�iQ��d�]�ʧO;_pO����N�a1�   ]��;   �U$��!�N��t��쬓ێ�Վ	����*��H����u�&���ct�Xi��4���n�]�k����ֱ�e�Ɣ�5/{�$iejJ�����}�:��ojuz�8!  �$չ9=��w�)��J��ggǊŢ*��fff��8+���[�0Q>}Z�׻]=F\�͒���    �VQp  @��eIc�!�N��t���%�p`��ϟN�5<<��׀��S����V����u2cc~�s5|��ٿ_��;hlEr`@{^�)�s��7�����&��=իU�  �Z�\��տRuqQ#�|�u�R�\��Ғu'��d�NU����`��cd�|X�  Ѕ(�  ���g�$�N�*;^p�Z8Y=�k||\���5`�p�:���Y��
��>U��W�^�b���e�����Sn�>����Z�����{��Wt���V�\��  �4z��[^j�������yӡC����f�9Q�O�d�ӧ�#�s�pϔ�����    �VPp  @7z����!�N�rt�p��-�=�e�X,���q��ߒ�Gg(��Eܯ �o�v�s���w��{�X��Y�lV{_�R�}�KU^\�ѯ]���ou�[�R�R��  ڬQ��я~T�rY#�z�u�9��jbbB�Z�:�S\.�W(�3�����;   �w   t_���C ����T�'��٬�0l��z����qEQ���Fg��v��\Nչ9�(#=<�}�߯=/y��{�Z�qN��蚗�L׼�eZ��ב�~U��E�z�!�h  ��=�;�#?��+^a�fG�(����>�F�a�a�h���=F\��$�H��k   �,
�   �6o�t�u�Ӹ:���p��U醆���yr����?��_��uS��k����u<���H~,f	Z��~�����������:��/�����U�� ��F��G�R��[�ّT*���A�<y�:�3"��SS��%	���z�n�4�F�  �E�k   �ē�/�C ���Bruf�:��VL���r���M^t���w[G0��M>����E���_�﹇r{���ޭ[��n�����;?�q�~��yֱ  @�5�U=�h��ǭ��X�PP�ug��i���][YQme�:�)���\��\   ���w   t�_�t�u��Zpwy��x�'�'�I���4�9���o�]A6����u��z�st�/��F��GI����P��G��G����:����jkk��  @�Ԗ����ާg�ɟ(��q�����������
�=j�DyjJ�]��c�J�RZZZ��t��[ҽ�!   ��`�;   ���e �T.���*ss�1̄�BӞ+���S�u�*�u�u���|_c/x�^������4z���w���ݺ��]?��/��w�[�R�:  h��c���>�z�leG|��������c�5���nRqx�YLp.�nI϶   lw   t�WHz�u�S�Xp��ΪQ�Y�0�MyJ(�}�u��	3������/}I/��AO{�u$4Y��_7=�����t��>��޽֑  @�?��&�����c�\�>Q�>3w���)��\<Nl���)�   @ǣ�  �n�A� @'sq�:;k�T�I��CCCL6s\��X:m���Tj����/��y��CC֑�b�(�u<�������Wv��H  �Ɏ�ٟi�ߴ��c�dR###�1z��ܫ���̹x�؂���T�   ��Pp  @7x����!�N�bA����m3&�
���7!��E*�y�u��	������^���݊g�֑�f��k�=���������շ{�u$  �,�����Tun�:Ɏ�r9��y�=��{��i��(�W�K��   ��Pp  @7��Z�:�e��p�r��}};z�T*����&%B�+�}�u���P�=��^������_�B�:�m�?�Y=�#Qfl�:  h���I=���Y�h���!�{l'�N�t����%g�x�آ_���   �h�  ��n�t�u����q��{荒��̄���m���05>>.oρޒ߿_�n�	����/�+>�y���)�p�����y�����}N���*�D @כ�����/}�:Ǝy����Q�ah�'EM���[U(�Sp�.��A�   ���׀   @���x�
\���*�ܷ��}���+�51���H(��u�-)�t��������Uzh�::\,�t�ޠ���E����s��0  zɁO|�'�TA���1'OZo�0�������̌ԇ�zL    IDAThX�0E�ؔ7IbR    :GK   ���Hz�:���8u�	*33�̄�¶�wxxX�D��i�+��:¦$K%����?�c�n��:�L<��m�����g4��gY�  �T�������u��H&����{<O�N�f�JE����(�����~�   ��Pp  @'��$�i���E����m.����+��59zEᮻ��f�0�Ϳ�Kz�_���{�&pcG
7ܠ{>�)��ۿ�;   ЕN~�˚���c4E>��Z����nW�v��ce�6����u   �RX	  @���:�@7pu�{��{��E�x<�!J���X2��^`�����O�T���
�����}������K�����4 @�i4t����$M�n[���̸��D�؂~I�   \
�6   �T���t����KK�1�lu
],����|ʛ���}�YG�@�H��w�[�~�����g=����=�� �u~XS_��u���}_ccc��b�Qz�vN�k�O[G0��2`�+)�   <+�   �DiIo�t�*���L����?22�(b�
W���d��1$I#��������6�g<C/���U���݊�; ��q��_�z�:FSDQ���a�=��	�.�z'���!�MÒ�d   x2V  Љ�!ik�M�a..ڕ���#����b������A/��P/~�i�0���?����~O��,p����u�g>��7X�  ��|�N���e�i�٬
Oo&�'��~���a�}@�g   8_`    x_�;�C ���E��ܜu3��+��6��d2�R���D�5���Ӊ�����t=��U�����g�_{����?���G��?�鞙
�S<O���.��y
2�s_��"����l��<n��L�;F}}jl3j}uU�J��ժ��˗����Ը�k�����瞻\^�ZM��e��PuaA�T=���%5j�m���p���Hw�}���n688���U-_��	lN�p��B��:�m���
I_�   �E�   ��%�t�*o������q>�i||��"���ݦh`@婩�����io~�����\�\
��z��ަ�3��o��Z�������>�ɤbɤb����>�R��K"!?����ףH^ɏ��G�bg�K&��bɤ�)H�%�?�5���cv���r|�R9W�_ZR��X/�k�Xߨ�U]^V�ZU}mM�rY��5�VVT[ZRuiI���WWU]XPmy����T1 Zm��?���������Q���<��������q�ҶEŢu3�܃ PE*�wb ����(�  ��Pp  @�y�u ��Ppw�f'Ѝ��)�D���t�:�g֖�K��j�G?��-������~�s���~V��o�����i���(Z/����TJA*%�l9�LQ=�J)�ɜ�?�T��l|��:���V�����ᗗU]\T}ee��_[YQua��}g����������_0� ��؟�y��%)C�������jp�ж}}��P�K���ʎܥ�]�(�[�_��%}�:    Qp  @g�Wҭ�!�n�L&�#����(���c�N�ې��t�}m)���ɟ�s>�!��b��LFw��oi�����ߩցE?�d�뗾���K%E���)<�1���(���s�Hn�=�����6��g�W��U[X��ku~~��kezZ�z�	" �b������J��m�iR��t��)�(�����Zsp'�z���ҒbH�R�����t�J��   �D�   ��_Z �����Y�f�6�=�N���6�h���oVr�.�<�DK�ߋ�t�;ޡ�|�%���u<���7�����k���Q�0�W��)�f�f7
�a.w��~�%�f�..����Ri[�ۨV7J��'���T��UuvV�UgfT��Uev���@7k4t��7]��X'i���-//kii�:JW
'�������]<^4�+$]'�1�     w   t��Kz�u���`���+�c��FGGۘ=��Tz�Ku�S�j�S��y��i�9�i�s�P����g>�o��o����}��٬���KNS?{��D�h`@�6�)�����BA��ɁOvvR|uaA�)�O��������˧OK�F�� ��䗿���z��X�:JS�������V��Q�N��zIezZ�]��c�q�x���Hz�u   ��;   :ůk��)�-J$����	�����ollLA�G}4���_����4��W�����+��i�@'��@��A���O��|E���m���
��(��W��+*d��ql�٩�Q��Ծ}W}|�\ޘ�^��Y�?;����*�:����zI~zZ��5��6�) wU��5�侮�u��:{2��Ç��t��������LQp����>$�u   ��Uo   t�QIX� ��kv��U�VV�c����b����[���cc��z�����<��?�sz֯��baؔ������b��P^,&?��?֧��7a��o{����5:v��V'�Q���⃃Wp��^|?}z}���*gJ�k�N�r�}���ևzԩ���+�KR:�V�X�����"��#��Pp�� t����H���A   �6
�   ���t+��\��.]���L&Ub"6Z`��/�q���}���w�lR*`�/��-�_�����/����g�9rD�J�����ߘ5��e�MN�2=�^�?[�?{����ɓ�-/�!8�]����+�=xbe�T���V>�{����T)�[G ��/K�-Ik�A   �.
�   ����F�@�
�@a.�_Ief�:���I��|���証�&
�2p�=:�����wM�I������_��d��Xl��~��~������H$�w�^=��Ze�2�&��RJ��+��{��Ֆ��v��&'U>uJk'N�=S�/�:��	�pOuqQ���=9���<���jbbB�Z�:NW��.h.Xs���H$�# ݬ��u�?4�   �Qp  ���K�t+�\.����'�>22�(������_�r������&�E���P�Z�=�������"{��}��@{���ѣG���h�#b�R��)�o�eS_[[/�OM]X�?qBk�N�|fR|�^ocr��N��=Yp��(�4<<��G�ZG�
.�+�ܙ��دI����u   ���;   ���: ��\\�sy�{�������f�Fi���W�Z���/����3s��酟��2��-L���y��ϻ�Qj�ŬSn����ɓ'5��W :��+�{���w_�1�jUk�Ni��������Z=s}��q�?�z�������~�[�Z*��jqqQsss�Q:^��ȏ"'�Qpw��dO�t����   7Qp  �����AR ���b�����sQihh�0\�ڷO��P����M=~���O���������й<O~�+�?�k�ۇ$=����b������� ��xA��Ȉ##�}Lezz��~���z���W��ۘ����ǵz����QZfxxX���Z[[����<OQ���'���]muU���<v$�y�h�!
�   0�۫I   �t� t;�*����Dg&�{����1��o�����w��׿.��W|�ೞ�~�
S�6%�	�[/�G����*�J�}_����Q �)�BAa����o���������ǎi�����ǵz��V�U�I�h���~W#=\p�}_ccc���P�*��]:Zp��ON���Y�0��13��t���   ���   +O�t�u�۹�X����L�}ppP�D�8\���������_��e3��^𻿫X<��dh	��(�o�ϟ�N�}ӊŢ|��	GU �K����Z������W�v�V���ѣZ;vl���v����r������?j��c�T<W�T�ɓ'��t����\S��V��;���$�_�[��   �=�F  ��$1z�!K�.ܣbQ�LF��ag���N�����%�Q������W,��a[<O^�?;�=�֯����P�<�=#����}?~\�F�: �	2Oy��Oy�%���k���.e����`B5�h�ᇭ#�E�P��⢖����t����Е�i�f(�M�:I�R���P   `��;   ,Hz�u��R)�mW����`&Q,jdd�:d2���#�����>=�#��%��xA�1}��;S��.����}=z��; \F��*��*s��W_[��#Zy≍��#Z}�	��<I���z�*��
��������8�Z�f�#�Ţu3e
� v.!��~�:   ��J   ,�O+@�6�����z�l��ص�*��
C��P��~��}����]w߭���<�MY���¾Q^���R;��t���>���Qr�m��q���V�k���z��>����������'$���j4���#���o��� ��Ȉ�9b�#9=���]�(�M�+�>.�j   �`U   �J�%�@�p�����lZRq����y�����)��뎏}�u;��Fyݏ�/(��w�����Ȉ�;f z�EJ]s�R�\s�}�J����Oh��!-OL�<9i����9Qp���g�r9���YG�8�������̸v�h�QI?/�O��   ��  �n��4l��M����ZG0H��}���9�0�s��5��B�<�wn�y���(���=%�˩�h�����Q ���a��޽J��{�}��e-OLh��!-<��C��/�;�kT�Y>x�:B[kyyY�J�:JG��E�f\���0���<�w   ��c   h�wY zI*����VUGf����X�:
�d2�ݻwK��VR����x���x|��~f������M���U��u��I�( �X*���nR�M7]xG���cǴ<1qA�}��AgO��f+����}����СC�Q:J,�V,Wmm�:J�U���#�J&�܁�M��$}�:   �@�   ��<Iϴ�׶[.;Xp��XG6���K�����Z9|���%xaxa���WNT�Y�BA�ZMSSS�Q  ��}%�ǕW��;/��:7�>�}bBˇ�����ѣj�jF�q%�R��ԉ��TJ�bQ�O����Q�|^�'�c�]uiI��5��u�DB����1�^�^I�`   n��  �vz�u ��$�I�m����PR��u
�0E�������g�Q��޽Zy�	�WW���g�:T����J%�j5�8x t� �S��[���n�W*Z}�	�LLh�l~bB+����d��T[^VyfFQ�`��J��������	�y�����>�=>2bÄk�!�6�YIC�؎   -G�   �2 �~�@�qm�Υ��'�p��w؊�bڵk����CI^(�g��N�Pun� ]x����ϿD�S�@�CCC�T*Z\\�� �&?�ڷO�}�T|�}�S��|�\�h��Ǵt� ��6*�<�\���<���jbbB�F�:NG��y�f��S��u��D��!���A   ��(�  �]�+ɭ&.��-��ly�rZ_1:��;�x��]�v)���?���U%��ډR��Ƅ��E�b�x\�3Ev/��Ȏ��<Occc:t�V]�	 z\T*)*����ܾz��z���ǵ��c��P�\6Jڻ�&'���F�m�H$T*�499i�#�ܫx2�v>��-�>*�j   ���;   �!��F�@/rm�Ε�{\R�I�Qp�����M��	s9��N�Tu~���v(�(�����Tv�����A��k׮]���P�R�� h��Ȉ##*�qǹ�u�9r�����Zz�q�>�F��v�O���`�X,jqqQ����Q̹\pwi7�'s��&��^)�ϭ�   ��Qp  @;���1�@/J$����EY_RAғgESp����A�r�-}�J����ϫ|�j�eϓE��0��<I%�z�  ��Wr�n%w�^�⍛땊V&&�|�}T�h�Ǵz��h����FFFt��A��_���u3���v�h�_w   �w   ��;� ���<�&Q���T[]���rY]��z�Tjw8���_�bq��K��ܳG��e���U[\ly������<�ɧ� �)�kllLO<�u @��P��W���Uz�K6n�--i���/?��}Tˏ=f�a�����Z,�"�J%�tx��$E���̸0,�r\:n��~I�H��u   �.
�   h�[%=�:Ћ⎕6�ss�Z..)s�����vJ$j�s�R)%S)5�UU��U[\\/]���E�bg�쉄b����C]�~�LF����� �p�tZ�[nQ��[���hh��1-���Z~�1-��?��׿n�T�#�+
ZXXв�'?��u3.Op����{%��:   z�~   h��Ir����k�t�/�{���/L�S��I��V�b1�������>��
�PP�VSmeE����K��F��F�z�7���XL~��ϛ���bM�t������jqq�:
 ��x�ccJ��I/z�$�{�y��}�8��'��522���^�[G1��K���]�:���/H�5I�E  ����  �V�Kz�u�W%	�m���9I�e�s9�����kttTa�޼XLA&#e.�gA�^�<ϩ]*��y����QMLL�\.[� t����)��'�c����XG�Qi``@����QLxA���OOx���)WB�h����J��    �M��   \譒��!�^��"]//�F�.]�=s��@���q����\�t�N��Sn��b����ƚ�� �=��y�uS��B��ܱ����u�rY��e�&\x���   -��   Z���^�ڢt�G����JmJ�����X,Z� p�D"���a� �.���Z��u3�J�:B�8�K��'����u3���&R��u��]+��   �M�  �*wK��:��\+�W��#�DVRx��D���bAhdd�:�K��r��r�1  ]̋�w��)&�_ �"8�K��ܥ���J\;vy�u    �&
�   h�wX z�k�t�,����6�����gttT�X�:��VE�1  ],���'���h4�#t�b��D"a����~�fzuW��q��`�e�ƬC   ��Pp  @+�~P@���k��<I�3_�&*�Z�.+�J���1 \�����m�_  .�r�=��g���<���Q�`�Lef�:�	׎�FI�l   ���;   Z�]�X= Z̵)T��y�M�'i��x�b��Q�D"�'P ]!�L�ȿ �m���:�?��Б��s�-�|�:��^�Y�;�Y[  ��(�  ��<Io����)T�F��cCI�-<�	�h&B�g``�� `[������}vު���: ���x<.ߧ������C   ���i   ��rI{�C .p��V]XP�^���4y���Y��@���a���N�Y�^�y�FGG)�  ���r������y�����c�M�r�}f�:�	��{�u    �VB   �l�b p�S��4����zE�ض�h�d2���~� �!�"p� `������Pp��T*�\.g�-b��0��a��	�[�� c/���:   zw   4�.I/��"�JYGh��ܜu���I�j�8��ϴ14��y��me ��P(P� lImi�:�>O]��Аb��u���<��Nq���|I�  ��A�   ��I�u�.m��+����A���h���řb	t5��4<<̉* ��i4T]X�Na&��g���b�������j���1LPp����"�   ��  �,���Z� \�R��&�%$���}Q���(pX<W��&���H$T(�c  �@yjJ�r�:���/7%��)��Χ���j�]�*33�LPpڪ(��!   �(�  �Y^!i�u�%.-�U�|��'i�K���@3��q###L|zH�TbG �U�=j���6oxxX�����N�{`x�v�t��o�   ����G(   �No� �&�JYGh�n/��I
���Ӷ�$�|��}��x����!� �G����fEQ��;>Eܫ���]4vC=    IDAT��Z�   @���  �f�t�u�5.-�u�@Rv�R�@�b1�J%� Z �N����: ���^p�ZG�*�b��w�	.�Wff�#�p���!|I�b   ݏ�;   ���"��K|�W��1ڦ�����|T(4+
600�X,f@���v� ���9b�ܷ��<[�h���{�	
7H�@   v��;   ���� ׸�8׭����νsy��E���=-�"8!
 p����Q���N�,�J)��Y�h	�O"w���H$�# .��S�!   ��(�  `��t�u�5�T�:B�4*U���clYLR�',��,p�����(� �ӨV���c�1̄ehh�'w�
��������XG0�ڐ����u    t7
�   �)R\�>խƲj·���؁t:�L&c@���R�d �a�T�\��a&>8h�k�b��|oᅡ����[���w�̽�ƬC   �{Qp  �N�%��:�"�
���y�[IJ7�y<�W����ع��!� �(��)�[�  t����:�������Z>���rp�ߌ�ֺ��w���&&��!   н(�  `'�,��V��.���\7��%5c�� ��׃[£=(���<�''� �o���:���޽��^/�4:Zp��˪-/[�h;����Ԝä   pw   �ă� W��8�m���fU��|�I�XG `���ϩ�	 �+s}�{r��]/�L*��Y�h*W�T�����v�7L�t�u   t'
�   خ�$=�:�*��*]Tp�%5s�?*��lpI��(���S� �Ԩմ���1LQpo���A�zhw1��ڎ�� so�   ��D�   ��v� ��\*�w����f.���b���<OE~v �e2%�I�  c�?��j++�1�x������1zB=�C�����w��^!��_�   �6
�   ؎P��Z� \����n)���2M~Έ�2���� $�� ����:������ ���3��|��r��{��Tff�#�]���],!�u�!   �}(�  `;^%�w�6]ȥŹJ���%yM~�0�o�3��1��Y�t�i� �y���={�#���4<<l�)\��^qp�{<��S� ���:    ���   �o� �.�HXGh��u��Ji}Q�E�B��,��*C� :'� ���=��u
S�k����sR���٬u����������lI7Y�   @w��  �����! ׹Tp��	�֧��BH1[T� ����sj� �9��:7g�T�O��Г�~�����&\:�t�7[   @w��   ��VI���9�0�h����>I�=7ܱ�tڝ� 6-��[G  �����#���F�=)î�%�O&�;:���	�C�р��:��0*   zw   l�� �3�Xk++j�j�1.+�z��e�O)[��v ���߯ �c  �l������LF��1�=�P((�򂸫S�]-��r�pC�~�:   �w   lų%��3�\�<U����pE9I^�?��xh�x<�L&c@�<O��� �Y��f��]��27�(y����6��U*��c숫�z����u��K&�� �{�u    t
�   ؊_� `�+����u�ˊ$�Z��A&����:����|>/�� 8c��U���R�y*�Z-��*�j���
-�KR�Ç	�܁��RIlY	  �M��  �͊$��u �\)�wr)��K�!�elR,S6�����A��	 p����e�\���#8app�:¶�:�]����Z���h@�Kz�:   �w   l�+�d�c��0W]X��pII��ƴRT,���+�٬|�C< ���� �f��;��$�Lv�ItA.g�w �^o    ݁�O   l����\'Np������9��Ci�f�R)��>= `�:7��G��a*�d����R�$��cl������z���C   ��Qp  �f�%��:�s\)�u������
mxt�d2�B=�M�9<� \1��H��uS}�x�<v8j�(�T��ϯ.�;q�@��r�"o�   ����   lƃ�X :DE�Y��m�}I��|=*��J�fLo����]9a �y����us�g>�:�s�Ŭcl���;���t��h}�L   ��hD   `�^k �9.-�u�����A�	����Ͷ� � �����: �Eժ����c���z�u�������[B��-.K��nIwX�   @g��  ���V�m�! ��ҶʕZt$e��z�q5�l֙� 4O.���  h���}O��y���(R��7[�pR>�����>y�~�r��w�#��:    :����  �o����Ң\'Mpϩ���Ƌ�6����lG:�V�1  -p�k_��`.s�M��:��<�S�T���i��)p�ĿN&�..K���J�3�   �v�   p5�� �B�,�5�..Z����Ғj�k2�W�ŔJ���@/�<O�L;�$ ���o|�:���3�i�i}}}J���16-�﷎`�2;k��9�t���WX�   @�bT   ��NI�Y� p!W媋�R�nC��jK�������[d�Yy^;� �K�٬f,6�}�kk����Q�����F��ڙ���S]Z�j5�VWU/�ըTT_]U�V[���8�=��j\�}au~�ү���z�r��jU���n�|_�M���Ӓnf��HlL���w�O$��E���|��'���XL�TJ^*�Lʏ��G��dR��� 6k��?�ڱc�1�eo��:��u��A���j��^.���*ߑ�K�;�Ҁ.�FIa   ���;   ��M� \̕E����-�������%(�2�٬u ],�J)U�U�(���yՖ�U[YY�,.���������UՖ�T]\\����������WW;�=\/����%�dRA_�z	>�T,�T�ͮ��I�����s��׷~�d6���z��׾f���Sp� �DB}}}Z8sBS's��.���9r|Ir�XЅ^"� i�:   :w   \N(駭C �X<��J���,��GŢ���[A�d2i@�<O}}}������&iT���ϫ�������/.RH�`��%Ֆ���\�t���{,�Q������\N��K��)��W�Iu]c����:����7���s���Z\\T�Ѱ�rEA��g���)���6܁�Jz���d   ���;   .��hXȕE�N([�����n��S�pu�lVSX�P6���ޡ�kk��Ϊ:7�����+����Ϊ<=��쬪�����ʊult��e��-~�����lVA.���� �߯h`@a>��XTX,**��L�7�|�{�:����>�:Έ�H�lVsss�Q���	��9��C��+�Ҁ.�ZQp  �%Pp  ���: �Kse�{͸���fz���bp�L�:��L&��T�լ����ښ*�O�<5����*33�3������(���4�����M����{�TRp� l��bq�v��M3��k�#Pp�,�RI���=���{'h'
�@G�]�.IOX  @g��  �KIH��:�KseQ�b�ؚ�݇f��qe��+�ri��V�<O�L��'�v�z}��>=��S�T��^/��>�q��}��%�@���������W|��)��
���B���RI��!Ň���b�6��ө�|�:��X*��ӟn�	�P�|^����Q.+�Y��n���{�0������u �%�^�Ǭ�   ��Pp  ���J�a��J��r��/)k��Z�f	\B:��ǤS M�N�)�?Y�����*�:��SZ=yr����e��̌��i�j���?������(VbhHQ������
K���Ţ<�o_��|�����a.w�m��=;�������:v��O.�8�0�Hhyy�:�K�yQp  ��p�   ���  ./�[Gh���kg$YΈ^dǕ��i� zH&��9���5�MN�|��N�\/�NNjmrRk�N�|�ʧO�Q�ZGp�z}����.�	�E������z48��X�z�DA����?���p	�XL�|^SSS�Q.)���/4�Q�ε	�w��=C�S%��:   :w   <Y��Y� py�Lp7Zl������q9��Q�V,S"����u���׵65���ǵv��N�\�z�V���䤓E.��ju��~��K>Ə"Ň��W|tT���.A��Ϛ��.I��ޱ�Ţfff:r���
�IU,=�:�@G{��Y�   @��  �'{���u ��ʂ�����K��K���
��:���d���^[^�(���8�ճ׏_/�ON2y���e�>��Ç/y��^T~O���tޒ����	��##J]s�u\����ɓ'��\R��9Ypw��?W��]�բ�  ��t��8   X�y�  �̕���|�_3&)��W��q)�t'�t�5�LFSSS�1�z]�'Oj��Q�=�գG�r�V�\���Z'����Zx�-<���w�����e�3��]J�ޭ��݊%m�L���a򺝦p��p������V�R��r� ������v�\��r<�b�Jz���Y  @g��  ��$�*t8�����N��.1��F�@+$	���z���ת..n�W���c����U��� HZ?	��1�;vɻ��A����(�'��Ur�n%FG��b-�t�o��5��e�w�eWqv���,�٬u��U�������Q�ƅ�i@xP�  pw   ��%��! \�rՅ��h�kv��vI
���KHM��<�S2����RS��:?�QZ_��$v �E��I�''5��p��^(>4�>�}|\�k�Q��k�SbtT�m���w��r'��a,�L���϶��M��r:}����u����u3��yE��u���;T����Iz���  @G��  ���: ��s��^[\l�kf%m�^�<^,� ������k��O ��J��^.k��!�>|Qy}��	5�����ѨV7~G�~���K��ܳG�k�U�k�ڷO�}��T�}���U��J�s�+?��c`<�S�X�)�1G'�KRev֩�;'�]aD�]��n   �(�  �qI�[� pu.L������Q����w4����x ��J�.��:?���t��F9s��-OLH�z�C@��--i�G���#��vm�Sg.ɽ{���$�����_��A��S|��#`r�����T�T��l.�W��#���Ӏ�zQp  �(�  ���J�C �:&�W��z�2�]���~��@�*��N5�u���[Y��?�C-:��C��|�ꫫ�� �I�Je���4u��dRɽ{�ڷO�T[^�	�A<�W��;�c`�Nq?q�u�wg�p<�?-��8�  �q�  p�+� ��0���.J���;iz�tf�;�$Lp�m��ꕊ����emM�3�������5����g�N��8����Nw�����H��D��L��.˒l˒�<�|���T���}�d��̋d�T���IR�7��U7sS�Ln���)O%�;q2�܉�+o���"%R�A �z��}_ �H �s��~��
��ϏZ�������2 p'�ZM�o��ŷ�6%1��Snd�tl��ࠦ��3�=[���`Lkv�t�X1�H�ݒ>-����   �,
�   ����N�`c�L�j�XpO��vI�����	�@�\�t )��
uE+��FC
7|���q
� �Ty�9��I���ww�rM���E�  �y�   I�&���Ѐ\Y��k�{Ҧ�KLp��\�����Ⱦ�����bB  zo��J����	�ss�#Ċsk U�"������\   �w   H�WM �9�,��Up�W���KR@��6ꀻV����{�l�Ⱦ������1 �ґ#*NL���mJ�w�X���*L@�>nm
� �k���%���    0��;   �I:i:��qe1�C�ݗ���W�:&���(���"u�u���
�uE�vl/?x�2����y  �m��ϛ��J���5��Mǈ]{~�t�X�rM���E�  �i��    0��Z�yHW��qLpO��vI�����a�[�VS��-�>��ٳjMM���k�]��|^����  l��sϙ���1�=	�J�t#Z�Mpw�`�WD�	  �i�  �WM �y�]�==~R��KLpǭ2��r��� �,
C��_W���K�ׯ�^h_��=���  ������Q�1�����f��c(;0`:��ZMQ&�ǥX,�� `k�Jz�t   �C�  �m�$=b:��se�T��I��.1����r�d��_+����P͙UϜQ������H���n�  ����ϛ��.I�wW�Ԛ�5!6�\S,�    s(�  ���Zd %\�6E���jώ�K*���;����X�+�6 ֋���gΨy�j"����B� ��?�Y��E���
��h������#Ć�k �����)  @�Qp  pۯ� `k\�6.-Iaس㗕�a&��f�\�t ;6��;�ƕ+�-��001a:  wT<p@}��o:�(��hxx�h���	��$ܨ�'M�   �I^�  @o�Hz�t [�B����سc{��{v����ey٬�H�,�= �֜�R���j��lJ�ؘ�a8  �v����聡�!���M&].�7ggMG�M�w �-_3    fPp  p��&�+�@ʸ0m����Oo4	C�H���Q��y5�]���t�M��yOP �N��������4h�|8�T���i�&�Kn� ,���    0#���   譯� `�\X��������ד#wOvh�t$w }�fSճg{��Y������  ���x@��q�1�#����<3K�.OpoQp�|�>a:   �G�  �M}��6���r9�z���Г���m+(��f�L��Ӂ�	�ΝS�l���me
� �����K�#��� Ѐ��y��	�T.\W,�5�   ?
�   n�I�! l���z5�'G��-ّ<�lV�L�t ��Zno�MG�&� �(������c��FFF������o�kw���z�t    ���3u   ���  �ǅ��v
�EIi���w�,�͚� `��v[���u:���Xy�>�  ��࣏*;<l:z,�˩����陌����_7:�������  �xQp  pON��C ��R�E�=��%&��V܁t��H��Z��tEit�t  n�祗LG@LFFF��n00`�uMkQp�_3    ��  ���$��bX����n��+i@�7�}�t �иrEa�f:F���� �0^���g�51)
*�˱�n�т�k�]X�+�    ^�  ��U� l�q�./��ez�$e��LG@�Pp��������]E� �4#�<#�T2121�=�Tb�$[-�����qap`�OI�g:   �C�  �-I/�`�\(�w���v���b׎�{�.�cm܁d�:�/]2��(� �f��/������e
�X_��	�R�$w �<I�t   ć�;  �[>#i�� �/�^���];V���KR�R!nB�H��Ԕ�v�t��˖J��� ������x�t�w��{gq�t��PpR�WM   @|(�  �嫦 �&�o�/)m���i�䣗(���Zj]�n:F��.x �e��?//�5���+����;��4�݅�j�垒�	+  �#(�  ��� ؾL&c�B\X�+l��r���LW��LF�B܄�;�\��i)�L��<;�  b��/�� C2�����b{=�'��Tpg�;�zYI_2   ��  ���%�c:���f��dRU�޲v����H��ʑ����Ph�M(����j�Κ��SLp $A���?���0hhhH��rv���?��y�bc���_1    ��  ���� `g\�2���԰���U���C���?��    IDAT*r ؚ���VOo�$߁� ��}��`��y��t���j�6�.\[�I��   �=VJ  ����@ʹ0e�[���]9J����1��� �Q��w�y٬�  �y٬�����H����X^'�K�>p���Ұ�4��X�"�i�!   �{�  �0$�� vƅE�n���x+����6
�@���u:�c����Mu �d��g�2	���T.�{�:^���M~��Я�   �ޣ�  ��_���
`�:](��u�w܌r;�L�9�b�j� ����b:ddd$��	�Ӹ�ε��MG���#����    �=
�   nx�t  ;��"\k��@R�;Qb�4	B�H���T�Z5#� &�����c����)�˱����������nziQ(LG �G$�k:   z��;  ��IϚ`�ྱ>Ii�3�7��$�+��%
�  �F_~Y�X�ĭ���z�>ܭ����!�t    �W�   ��yI�! ����¶֓T�^��Qp��(�	Ej9Tp�)�  L�d���_6�	T�T��~O_#p��ީV�(2#.\[�   �Qp  ��WL �.L��,-m�gKJ�I��� ��jUQ�e:  �|���7	�y�{����Ga��w�K
�U�4b:   z'�k�   ؜ϛ �;\X�����/C6��G"G��i����Oi�i6MG  8j��WLG@��t�+W��ήǤ��# �x�^6   �C�  �n�J:d:��pan��
���F�]v`�t$w Y\)��2� `@P�h��L�@�e�Y������A��t��y�b����1_4    �C�  �n_1 @�����f����&0�7��$G�VS�n��+
�  �~�K���;344Գc�Lp�^�<*�E>+�7   ���  ��^4 @��>�=
Cu��-��/���8�����EQD�H���.�f�f�t ��F�l�\.���H�r�ݡ��.� 2$�1�!   ��  �U���� �����Ғ��BoYR��qb�0 ���#�,o�w @�*'N�t���H������傻K�ym��8��   ��  ������ ���	�-�LFR_����/��	�1�0Lp�[-������� �۾�~�t����<����.���m��8���  ,E�  �^_6 @w
v߳ҩն�3I~��Ď��XK��# �s��s����~ �9��A�<���H���߃2z�g�-�����^ۯ�zH�^�!   �}�  ��Y� t����3�ݖ��R1	��tLG �����lИ�3 ���_��<��w�}���]?f&���h���P����k��2�^6   �G�  �N�I7@wپ ��b�0���M��Lp�(��EѶv�Acv�t �C����H�R��|��W�L�O��C�^�w�8v4  �w   ;}�t  �g�ʝjuK����xd���5Pp���뒣�6��MG  8b��I�2)544��c��]��N��ҳZ��   �Pp  ��� �>�'��[(�g$�{%v�N�ÝQp���W�h--)l�L�  8b�W�t�X�R���]=f�����Eۡ����� GHz�t   tw   ��Iz�t �g��V��E�uB�4	D�0�Ղ{cv�t �#���y�Y�1�b��i``���tv�{����4#Lp����    �.��    X��$��*
�#�T{qq�ϵm����y؁�;`VX���`w @\����<�o�F�v��qW�;S�)�����    ��t    t݋� ��'�o�H��}w�d)�c�s�fS���6��LG�+2���e�Y��2�//����+�y���ok�K%yA�L6+�PPf�go�����-�(Z���Y\���_�����ӑ�h�9�Z��V��Q�|#g������QX�)l��?�Z��X%���W�b:,P(T(T�׻r<��{vd�t����X�I{$M�  ���  `�gM ���å�M=���&ܱ��7����te��+�# ��\N~_�����r����������BA^���_�>��+��W(0��&a����T�h�S��������ZM�jU�jU����U���:ժڋ��ϻ���u�UE������'�Pq|�tXbppPW���	�����ఌ�/J���   @�Pp  �˸��M� �}��)�͚��S�ju��d$�z%vܱ
�9����˗MG@��~eT*
*eW>n�:�￥���SJ�o�F�n	�M���o�h��������:��˓恘��Ϳi:,R�T499�0w|�`e��Rpg�;`�E�  ��  ���� ,��t��&&�$����l�b:��j)�"e2��ĭS���`��ŋ�#`�2e���RnxX��e��)�k�G�������y�S���\N�]��۵kK?�ᭅ��Y5�_WkzZ���պ~]͙�ffV��:��.`��'�������x����>�����X.߀N�����Yd:   v��;  �]>o: �ޠ�������X_Ej����� $N)l4L�0�	���J��ݻ\T޳g��Ȉ���˟W�칡!
�芌�);8��ࠊ���E��쬚��j_��\���QsjJ��5�^UsfFQ����H�L��o�������`w
�Lp�w�j{$=(闦�   `�(�  �##�i�! �F�P0���Z����Mm�&`�;��j�(�1[-)M�0�	��V'l��Wn�.eW���޽��ݻM�6tc���h�ϫ95��q횚SSj�|��u��e��v�]_��J�����ee�Y�Z����])��0DpܗE�  �
�  ��a�! ��oQ��\(�����䱍W(ȳ��/�o�� [��#�i4T�~�t�T��[���ޭ��=���{�*72��
�.P00p�rs�n�53���+jMM�~��/�q���W��y�����1�F7���7�a:,V�T455��c}}�x�"o�q���w�z�����C   `�(�  ��K� �����S�!�	.O���(����Y�tI�"�1�+�Qn�.�Ɩ?��S���J�=��3�H�L,��gϺ�	�M5�\Q��U5�\Q}� ߼�k��,O*/�ױ��]y�Ns�QpW&#�TR{q�;�Rĕ����� �	-oz��B  �x�  ���  z�`y	�S������e+��`�Y@��f�tc�Ϟ5��LF�ݻ�߷O�����7�:?:ʮ+@x�����*������̌j/�~��.���~�W�*�tbLe2����}��1����r*�J�np�a#A?w�1��^A�3���A   �3�  ��'�� z���R��1�0!��7	F��������3��2��ܮ]�����R~ttu{~t�;`�����x�۾��j\���J��R|�]����j��Hl�������_4��J�]�/w)Qzt6���(�NxI�  R��;  �^��Í��ŷ;-�f$��;���t$X��TE�d2�� �p��~���;��r*�u�
���Qؿ���e��#0,�N�uך�o�ͩv��j~����?�����߷a�k_��7�a:���/�����N�����X�s�   `�(�  ؁�u��l_|����$/�(�su��E���
���(��VK
C�1�IK����?*���o��{�*����@����+�?��m�[-��(��;�ڹs��;��^7�6���������ۦc�1�穿�_����>���Nka����R��m�%�$阤]��L  ��Qp  �çM �[�/��iJX9�&�.�c�(�����i4�x����Ri��~s����r{����Q�ߣH�+WT��CUϞU��YUϝS��Y5''̈́5(��:����~��LG��*�ʎ
�.����2��8���iy0��m:   ���;  @��H��t ���w_�ݿs�α9�F�t�a�e:�1�g�(�yz}��US��A�TqbBŉ	�&&��5 �H&�¾}*�ۧ����[�juy����k��-�9����~�������}���|��Q�R��\.��6o^ty���Ғ�� �y�B�wn�(�  �w  ������Q �����:܋�2�F�wl��;���׳c}}*8��]w�|��J��p�]*:$�	� ,�J�;vL}ǎ��xgiI�?\.�����+�K��(2�vg��zJG�w�۽�t@����������e���[�z�gl��d��f9�����    �
�   ����  z/�˙��S�uPK1�0���p؜Z�f:������;��� ��¾}��Z��^:t�i� ��\^��ޞ���������ϜQ{n�Pҍ���ա��w���LGVn��8\p��a�6�|��;`�#��K�`:   ���;  @�}�t  �g}�}�o ����|
��@��Q�ٴ�� 	\.�_{�M=�/�U��P��A�Tqbb�c|\N����8�ʉ�<ޜ�V��-����N����vN�PR)�T���_�]_��<�wC��r�m��=���ۋ��#����������t   lw  �t�/�� z�����&��0�]���~���j��;��т{kiIsgά~��<�GG����Tb/<�������r##ʍ�h��GW������������xs��!���]�/�,�P��k;Q�T499��sy��z;�����l V}N�  R��;  @�}QR�t �g{���;ܱ�ZM����c v�"E��F\��/����ݿ��*NL0� R����w������Ǣ0T����;�h����;j����J�k�����_P�}��4:���
�[�v��n�u6 ��1    �G�   ݞ3 @<�٬�=��؄��ʇ
�؄j��pX.*�L�0��/~!Ix�!��5� ��Sq|\��q����Wo\��\x?}Z�3gT�xQ͙�gg6��?�)74��ؘJG���{4p��r�v��-ۖ�fU*��|>�;\pwe����� ��t���L  ��Qp  H��M ��-�������h6�j��
.� ����vI�Z)�'&' �J~lL��1�<���(@��\p�
yA������X�EQp  H%�t    l�I�M� ��N��H�z���J����wlV�V3�Z�阎`D��h���$I��q�i   �k``@�Lf�?�\�2�������:��|�t    lw  ��z�t  �y�TX�*
�կ�|sqb���0���թ� ���	��o���ʟ/Lp  ��}_�����s�ft&��Г��~�   ���  �^�1 @|l�,��XiץiA��H�EG&���:�����_�$�TRnd�p  ��T*[��x�Rp��:���t��   �:
�   ����  �c�d��O3r���;:��l6�l6M� �����?��$�t��    =���'��ڲ���ێ�f�u6 k���    �:
�   �4!�� �c�d�v�����:Quu�۷��4=��(MG�]��u]�IRq|�p  ���<O�[�A�/�t��G:��R���s6_g��gM   �ֹ�   ��L /�'KuW]4��&�c�o��@w�Xp�������  �k��r�GI�-
C����=g�u6 kz�t    lw  �tz�t  �y�-\��:#�
�ف��2�jU��� #\,��������m0	  @o��ey���]�!����a6_g��QIGL�   ��Pp  H�'L /��N��p��{'�./�c{�0Tu� ����(u�G?Z�:O�  X��<�m�<pt��$u8��:�u}�t    l�k�   �t�t ��<oKS�Ҧ�Rpwmz�$[�"����� +�Vp����՘�]��	�  �v�[8w���^\4��(�Nz�t    l��	   {� )c:��ؾ�֩�$9Zpg�;�aaaAQ���Ǳ���?��[����e(	  @<���6=@���A6��t �{�t    lw  �����  �e}�}iIyI�� 0���n�Uu`�x nQ�c:Bl�0ԅ���[�  ���y*or2�_*�8Mr�(��~����K�0   �G�   }�4 @��٬�=�^Z����.O���,,,�� �ǡ����Ǫ��|�@&#���   �Կ��]�q�C����7    �G�   ]vI��t ���j*�a���ؙ��yE�qtׇ�����I���4   ����Wf�{�MNz��wۯ�Xw  ���  �.ϋ�p�sl�*���M�0����8��:���ժ��U\�i$l�u�/��Ǽ|�P  �xy��Ri�}䂾>go lSp`��M   ��Q�  H�O�  ~�/���u��	(�c���MG ��H��ʫ��17w�c� �K6|N���;�Ʌ	�� ��#Z�)   )@�   ]5 @�l/��].�;��9vn~~^a�� e��ɟ����   ���߯�&��}}1�I����=g��6 �ʈAR   �A�   =r�6@�l�*U��%N�lbj��0��t������Wu��Q�c   ���T*m�<GoJ�T��#����� l��   �9�  ��	I�! ���R�lVrt����st�st�����=(����w�i6o{<l��  0�o��]-�3���4    �C�   =>c:  3l�*U�Ė�����U��T��M� ���韮�xD�  8�����z�.-���s6_k��㒘:  ��  ��q� �a�T� 8\�6��lS�l���~��>X�{Lp  ��f��o��Z�h��S�[������ lJNҧL�   ��(�  �� G�:U���_�����Ip边�9�ah:�~��*r�O�d��E�v�I   ��o��r�T�)I�Da�N�j:FOQp����    �w  �t�W��! �a�[__��w&��[�0�����@�Y\p������}o��G��"n�  �٨���1%Iۯ�d�YyU	�aO�   ��q�  �L� fc���<�J%�L;�izzZ��[�ؾS���:����w  ��b�(�����O��jA�� ���$�{�;  �%(�  �Ó� 0'�˙��u�RI�穵�h:�1�nu��h6�Zr�� ����������w6|^�jŐ   92����Lx�Yہ�56� �iÒ�1   wF�   1 �96.��X@va"�z\���133c:�jK���韪1;����  \t�����y{ہ�5�|�t f=k:    ;  @���I�Ӭ.�;0l=.ou��XZZR�^7H/�Q����6�ܐ�;  pP__ߺ7:�<�݅�A�� �,vN  H8
�   ���$�t ��r9���P(���;ժ�4������S܁��x�]*��?��>�pS����  H��TZ�����v&��v����4    wfߪ  �}�2 �Y�Mp�y��6܁����W��2H''�����ݦ��N  ����3�����Ё�����'��?�  R��;  @�=b:  �l.��\�syz'�"MMM����m�/���z��M?�����4   ɵ^��+�{��Y.$��z�-���  @��yF  �.�M `�M�|�W�X\�څ��O�Co��ͩ�l����e�_~��[z>w  �\.�|>��LF����S����s�Hz�t    �ϮU   ����t f�Tp��T4����#Lq�Ǧ���}M��Ɩ~�����   �Mq�o�I�%mvܳ�z�m{�t    �ϞU   ;=c:  � 0�k>�`:0l=>w���ܜ���@�XRp��H��ַ��s� ������;��Z�@��	�(�    IDAT� $�0    �c�  �^O� �����N��/�<�=Xg:�-Lq�&���#t�����u�ԩ-�\k~�i   ҡX,*�������;���=�w ��I��t   ���;  @�}�t  ��2Q�P(��Xy���D��0��6??�w`l(�Ga�_~����Y&�  �y����鞫wvܳ�z�{�t    ���;  @r�0�y�,�ݶ�w�M�詫W��� �����ǚ{��m�lka��i   ���r�ܽ]�IQd:FO1��

�   	E�   ����  ��e����;����Ҙ��<y���p��Ғ(�����{kiI��ַ���m��   ���~�0Th��`�\o�c��   ��Qp  H�'L �6Lp�<O���]��z=^����)9�199����{@7�����o}K���m�|gq��i   ҧP(���{B�����N�f:BOA`:�dxXt�   �7i   �u�t  �`C��X,��X��傻��T8�W�ͦfvPz\������z�?���	�   ��>��w�݆	� V�$3   ���  �\�M `��yVL����d�B靸�@3����n�M� -������N���c��_�R  ��*}�|�c���(����   �v�  �� �n�! �g��vI*�1���;��0u��5�1�dKi����K�W;>NkfF��.$  H��_��A=���n�@	 ]��    �w  �dzT��V ;bC�=����w��Pp�����:����L&#y�\�i4������+l6�^X�ʱ   �*���r�wx�{���G&���	�   p�t��   ��1� $��mkMo��.��O��Y�/_VĄf`]��Mq�[�����];^sj�k�  H���cx����_�����yP�:   $w  �d���  ���	��ܗ�bN�>�aH���V`]i*�_?uJ���v�����   �n�����N�f:BO�p�@�$�o:   nE�   �>a: �d�a�m݂���w�w�4==�F�a:�Hi)�������O��]=.�  �R��L&#����m����7    ���  �<%Iw� Ҿ]r>�W������wB�&EQ�˗/+�"�Q��IK�����5���]?nkf���  H��T($�}�n�`��_s�u��   �[Qp  H�G%�����O�*�aҙ��`���@\j���_�n:�8�un�J�����Ʒ�ݓc7��{r\  ��)���RIZ���ۯۤ����;a:    nE�   y3 @r�}�T���:KK1&I��	pH���I5�1�DIz�=�t���ծ�{r���TO�  �6��32����0�����~�@�= �;_   ��;  @�|�t  ɑ�iRw,�[����0�IE�.^��(�LG#��_~�ۚz�����;  ��R�����v�ћ�ۖ_�I�57 ]��r�   	A�   y2 @r�y�T6���b��[]߉���H�F��k׮��$����˵_�Bo����5���==>  @Zx�����v�X4��&�p;,  $H�G  �'/���ve2A�V�e:�5�<M�N��%��LpG�LOO�\.���@b'�7��o~SQ��uW����   iR.�U��8z���;�Qp߾ ���$)�ϯ�vpC��R�ӑ�|c=�"'L   �G��b  ����fEjy��Zn,�*
*
��.�*���r�ӫ|�_-_g�Yy��D�Z-�+E�z�.I�t:j6���j�������V�iaa�Y^p_Z�)I���0�.]��ÇW�W%�����O�t�R�_����������  @�W&���Np���$���r��*�����o�\*�n�6\(��n
�t:j�۷\���z����E���kiiIQu�wl�æ   �#��  $�I�`�r��J���h���k�w��r��b�V4���iaaAsss����������477�v��͸���Ŷ�/�މ�ۛ#���.]������<����i�Ip������_c{�������z]��Eu���K���j��+
C�u:
�UE���KK��m����v[�g�FC�7_F����d|_�:��bQ�lV^.'�PP���J˻"��;����LFA�,�X�W((��_*}���@�) ���q]�su���;����fy��J����!��Q�T�u�v�|ߗ�����T*>?��k�7_���������f��$e$qw  @��  �.�M@�y����!�ݻW�������e�$���ڳg���ٳ�����t��U���hfff��6M�I�b�f�:پPz'LpG-..jjjJ�v�20��	)�_?uJ?��ߋ�5�/�|�h���Ya���쬚ׯ�9=���Z��j�Ϊ15����G%����YZR�������岂����~e+���
�����GvhH��Aeؽ �5�(�w���NGQ����v'Y&�����X�^1��kddd�cϞ=ڽ{wjw��<O���\��KKK�����̌&''u��U]�~}u7Q`��%����    ��  �4��t	�@{�������E�RQ&�1-�rY���ÇWk6����ֵk�t��]�tI���S�LZ��M�].��:��w��5
������	i�I�qk�������R�^��u/_���$)
C�ffԸzU��I5o|�vM�+WԜ�Rsz�����j˓�gf���A�����j�=;<���!�FF�۵K�ݻ�۵K^�S> H���.*�jW��ZZp��w�Lc�=��ittT���Ӿ}��{��M]��I�\V�\�����c�v[��Ӻz��._���/j~~�`J��IQp  H�t6%   씑t��H�R����Q���illL{�����[�r��ŝ�~X�T�Vu��MNN�ҥK�x�bj��Zp/nb��咚��ߐ�.]���7܅�U&�Fa����h����_�ޣ�{{~^�T;~��~�W��95������bc�9��椳g7|n00�\x_)��w�Vn���Sᮻ��} �*�b����ZMZg���r]�\.�9���<�3+qn�ٻw�mׅ/]��K�.��ի��.c>%�L�    w  �$9*i�t$K>���Ą&&&��~U*ӑR�T*�2��nkrrRgϞչs�499�(��\[Z��f��"���ʣ8��t:�x�&&&X0��2٬�z�_�k]�����N
�Q��ڹsZ:sF�>P��2{�ɉVh�ϫ=?����4�*�o�
��}�yll�?6&߱� �ts}�{'�݄�M�{����y�������W��H���u�K�.��ٳ:{��f����	�   �,�M	   ;=b: �addD��������O��� X�x��O�V�����:����}---���*�w��������N����sx�ң^��ʕ+3��g���������?0���+W6~R�q��O�V��-�|��=��l�HkvV��Y-������Ua���SqbB��U�� @�����3Il/�'�ׄ�����5>>�g�yF�jU�Ν�|��gϪ�l���4    ˒s�  ���� t��!:tH�p�5��X,��ѣ:z����y]�zUgϞ��ӧ555e4[��6k3���ZI����H���9��y������*c��ޙw����M���2kMpoLNj�7�?�|S�o��N�j lpc
�ҩS�}���T:xPŉ	��U:tH��	'&�s� 0�oh�tcl�~c��������w��5a�J���;�cǎ)C]�xQ|���{�=-,,��3�$I�n:  ���ה   ��:���=�ܣ#G�(�˙���LF�����?���y����z뭷499{�4܋�غ������;RdrrRA�R����&��y�����7Sm�����f~�U�{o���0�n
�M-�:��5����{U��P�������*=��ࠁ�  ��)�[+��n��ittTG�ս�޻�kh���y:p��8�g�yF333z뭷���o'j�O�\Fҧ$}�t   ץ�)  `��M@oy������رc��Sd``@Ǐ����533�S�N�ԩS������m-�۾@z'LE�\�|YA���p�g��ުV����U�P$�"��w����mW��q��f_}����{��|���>��W}�ޫ�訡�  ���`L�^7����vs���ѣLjO���a=���zꩧt��e���{:u�ew7�w   ��ה   �Ӱ�}�C�7FGG����{�Q>�7;0<<��\�?���]��7�|S���=\�K[�=�ɨP(l��w 5�(�ŋu��An΂2�/y����^�n�~��u}��� 6v��>���XP����{�w�}˟�Sq|�`J @�����I���a���ܳ=��uxxX=����>&��\&���ؘ�����OZ�ϟ�o��3g�(���c�e  �HWS  �^'���!,���t��ꡇҞ={L�A�޽[�>��>��O�̙3z�7t��yEQ���I[�=�����׮VcH�L>��H�N��?�PLݟK�vx�\le�������~�k�h��i��Wo���V��	|��?����2�� 6���)'����lP��~׏w��=���:p��2�װ��y�����Ą��N�:��^{M��Ӧ����q   X�  H���;��ٳ:�������n1<;;�7�xCo����]*p��H�ىT�O �o�$j�Z:����ǻ^ �&��J1�]����t�?���� �53���}OS�����
�'Oj��1� �T~�L��Rݺ~;<<���_>��v6����z�!=��C����/�K����j�ۦ�a�J�n�  ��jJ   ����}A��������5<<l:��O?�'�|R�O����s]�|yGǴ��n���,t"����j�}3�5 i�e����5���?ԛ�����U ��������=�<��o|C�O~�t4 @�d|_�BA�ެY�{��u7��t��w�ĉ�b*�ў={���~VO=���x����kZ\\4�W�tD�{��   �,]M	   {��a
�J%=���:~�8�yp��V��ONN��^�;Ｃ0���[�LpҫV��l��y=މ����~�/�EO_���f_}U����ܮ]|�UyDC�>�<�5 ��b��?IӶ�����n�\N<��>��Oj``���f�BA'O�ԉ't��i���?�իWM���w   ��Ք   ��=�`�u��q=����+#~{���/���{L�����x��Z�M�|���}_�|~S��T�=N�\�&o �liiI.\����)��J��?���Y?�g��g��3ͩ)M�ٟi���L��w�F�W����J�� LɖJ
ff�6$f�(��u7��`+n�r��%��'?�|�(�LG��}R�wL�   pYz�   �: i�tll���:y�&&&(�a�*��>����G�믿��^{M�ZmßKS�}+�{�/�މ�"(,�����/ꮻ���EX���zr�����G��+�Ʈ. �X|�m�~�m}�/���|�K�C�]�L� �,(����+�o��U�m���ȈN�<�{�W��Ő
���/����)���?ջﾻ��>�M   p]z�   �:a: �l߾}z�'4>>n:
,P,��c��ĉ��/~����j4�>?M��&�w,_ ��	���.]����1J�J/&����?���?P��t�� z������G����j�k_Ӂ_�u�c b���Krm?����o�wx�?00�GyD<� �vtŮ]��/|AO<�~����7ߤ�l�L   p]z�   ���� Xۮ]��裏��ѣ���B�lV'O���?��_}ݢ��ڒ����xLp�e��������O���x�2A��ݝ�������D��@X��¿������#��[���K�# b�LpwMd�|����X�}�Q��虁�}����'?�I��G?�{ｧ(�L���I�KZ:   z��;  �y���[������=��CQ=���t��I=���z������L�fs��k-�%Ua�����;a�;l����?�P�  kd�ٮ�O}�;�����"&�Vi����o~S������{�i� `9�XTV�'ɥwu�(�y�D__�N�<��z(U��^���������)���ݓ������M  pw   ���0!*���z�)��0�P(�����?�W_}U�����0T��-��m)���w�wتZ������a/�U�ÿ����ٻ��8����OU7@c%A�$���H��(J�$j�D��,ْ'V<��ؙ$g�8v$'���M�Q6*���ڞ��3�=�NNb'�8�sm�VdǋƖ-J�@�;[�F7����H���4��~����spD��>�����~��?��SEJ��z����ڿ_�>�	�o�� *U4�#�J�囯��hT��պ馛�m�6��b��z��t��}�;���ӧmG�w   k�є   �\��5�C�]UU����z�p�\Āu�x\w�y��mۦ�|�;WL��Lo�4��`�E(������K������sc�Y?����ɟh��?_�D �j��i����?�#Ϳ��q  %��%���n�y�\NN@�Ö́1FMMM��_��/��lZ�d�}�Quuu�[������lG���v   �0c�  �]k%��V��hӦM��>�]�vQă�̛7O�x�;t��)��^]]=�Ǉy�{���v��FGGu��1e�Y�Q�9�m�'���{����ہ�ɧ�z�7S}����( �p/������)�TJ����ZZZ(��w�����Oh��݊���k�f�   �;  �]�l�ŋ��Gս���E����^}�U?~\����Lj��+��h�\&�#�٬�;�t:m;
0k���>64�o}��:���W	�;/�ӫ��[��mG Y��	�aSI��������K�x��F�s�N=��ڲe�Ǳ)���   fQ�   B��eV__��o�]�ׯ�(�1F===���W[[�.\h;�[̸�^AGg��;�"������jkkScc��8��ʹ�>|������h���%^6�W?�qm��C5mm��  ����*I�$c5MyUc�N�>���ny�g;P���z�}��ڸq���o����v��Y.�FR�  �  ��v��pG�6m��?N��5>>��Ǐ�������b4U4:���+i��LE.\���S�N����v`ƜhTr;}z��W�����r; IR��O���o��x& ��\<�w�	rAR�J���~�={�r;���M�}�{u�w��*�{IX�J�`;  @XQp  ���u477�]�z����O��hxxX���שS�d���a��w����_nLpG����̙3����D!S�_�����}������!��H�߯����ڎ (�H]ݥ_�l���ꐂ���<x�W�"��r]W۷o��?�+V؎&[m   ���`  �7kl�d��jǎ����Dl�����g�jppP+W�T�eZ˭��zfO0�"���-&�#���d�l�2��!0�Xlқ��|^/�ٟi�_���� &p���½{_��v �]~�zL҈�(e��a�t��	e�Y�Q��kjj�#�<��^{M��/�����v   ��b�;  �=K$5�Q�Z[[����G�w�܎�6::�����ֶY���|&�"��ʉr�9�+����ѣ	SA6��L����k��?ڟi ���r�ڷ�v @D/,��uM�
�\NG�ё#G(���9���7�}�{�֬a�R�m�    �(�  �ö�%ຮv�ڥ���=jmm�(c�zzz��+�hxx���ϸ�Э��!2ÿ+�]�&���� �r&(��߿_���:���[H h���]���� �9�|7��܃2����_��������(@����顇�<0�]6Q���   �w   {��Pi�s?��h�    IDAT�sڵk�\����l6���̙3e[3�(6�t�ɘo��^vA���n�:uJ�|�v`R�Op7���������?h��?k߉?�s�  s���o�ZR��f�|~��'N���K���� V�_�^�=�����lG�D��&  ��0{  ��ѦM�t�wθhTc�N�>���A�^���{f:�]b�;�7ittTmmm�_V��b�=�߯{�i����-'D����F_]�+Wڎ ���U7��$��J��{:��ѣG��qF�\. z饗��/��<ۑ*E��U��X�  :��  ��m� �����׽��K����Ȉ��߯�����3�}��.w�-r��^�uuww�c;p'Q�O~�������̞1:��/�N ���
�aፍَ��uww����ہ˸���;w��GUss��8���  ,��  `�Z��n���z�'�a��Q _�<OG��ѣGK6��	�3s�q o:���;�l6k;
 ������O5��c;������$n����\��T��6������t��A�8q�	��$/^�����\;)�km   ��� (�O��K{{{c��Ǘ8�s���3,I�H$��  ��^}�պ�~���l�*�q�}�v�v�mr]�����ק���Y�F�E.X3�}f��L-����ѣZ�h��`U&���ӧ566��+4��K�#��s�4�ӟ�q�V�Q  ��D�rc1yn�S�=�	�TJ]]]�𽋻�.[�L���7�!djkkw���A��  T*�q���|��u��ncL.�N���d?����Pp��|�3���������ht��yˍ1K�i�Ԩ7vȫr'b�qFFF.Z�1�n��I  J���0��bڳg�֯_o;
(cccz�״j�*͛7�h���|Sn�GFˍ�;0=��t��jɒ%��>̖1F���:����f��V��b���w 0���R�=r�#o5Qyx>�e���['O����6��mٲE---��W�����q������|���s  �߿دQ2���8�������4d�9�8��uO����D"?�����?��tY� (*
��L&WJz��ݒ6KZ�8Nc*���$�u/�q�8�[�ρ>  �r��9�i޼yz�����b;
H�穫�K���Z�lل�3��f���߶�.�78K������5��9���N�u��Y�]�s*N�@����jկ��� �Y���|��
I�����t��1���[�Y[[�{�1}��_Չ'l�	����ێ   .c�q��!YTR��&�q�K��y�\ו1F�TJ���9c̐���^�􂤿��'_��@�(��Ѕ2�c��q��Ƙ����� @p���؎8���ڻw����mG���[���jooW4:�����{���P�uwwkhhH�/f�D>�Woo����&�z|��2'P���Xw��[[mG ̂{��H��0��y'�ɨ��K����2 �"��Gы/���������Ȉ��Ƹ> @ c�$�\��,�QI�uvv�c�$��uIE��(��@2���u�_�<�m�VH��]1Ev  *Ooo����8�n���ܹ�ɭ@�R)���Z�f�����^#���ya.��55�# ���d���k���Z�`��v� &288���n���O���%K�VW����"1F�/���?l;	 `"W�?������&���ѣ�v10w��j���jii�?��?+��>sg�Qoo��.]j;
  (��[/|�)����䘤��~���>��?��ܭ���?�4�N��1�~I�$�80  \�ΰ0�HD{������mG*R6�Ձ�j�*͛7o�ϯ�eY;�A&��g�����500�h޼y���Y�d2:w������u\W�+Vh�С2$P����_)�@@]]p˅v�͖}���n�<y�Ap@�lܸQ����������!�={��;  ��Z�:���I��d2��t�q�����?�Ї>t�r��	�q�u����H��1枑��E��   ����mG���Z=��Cjkk��h�穫�KmmmZ�dɌ�;�	�&�A�	�����y�;wN���Z�hѬw�@8������G3z^|�*
� �����M^6+w�� �\}�:�K�ĉ���.�@-Y�D?��?�/}�K�����zzzlG   �����ydd�����!c̿������Ǿf;\Pp/�g�}vw.��ϒn7�0�  HzcZ$1���ܬ�~X��Ͷ� �q��i�r9-_����ȳ-��y��K�(�L&��_]���jmmUUUX�%�����ק���k6;)�W�.A* a�O�5������lG ����#�\I��Ow���x���G���fT ���ԤG}T_��u��I�q|����v  `�1�Q����ݟL&G%}�����>򑏼`;[���^d�>���l��v�\.�`;  �s�α�������C�����r�����ؘ֬Y#�u�|l,��1���<���m@�)�J���I,��+c400���^�����ujW�*^( �7��Pp� r'8���T��{٬d�T�@����r:|�0�a jjj��#���_��^{�5�q|��;  �J����\no2�Lc���~�#���l�$܋ �HD������p.�[V�C  Nl�:�M�6iϞ=�.�����!8p@k׮��$:��������ࠚ���p�BE���
3c������۫l6;�ף����C�  ��j������ƹ�R���d2:t�PQ޷��H$��{����Y����l�񥾾>�  �58��\.��d2�'������G"��Է"�J�ttt�$��u�[�1�y  @0Pp��Ν;u뭷�����^{�5�_�^���>f����;�R�XtRss�ZZZ(���1F�TJ===E-��W��\W򼢽&��J���##���َ ���$�0�g2%9��N�u�С9��8�Ѯ]�����o~�����N�5::���  `:�%}�����;::^���SO=�o�C�1g�����d2y�q��9�s�v  0lc�V;w���ݻ)�>��fu�����N�u
�C�(����ק#G��ܹs��r�#��<�S����t�ԩ�Otc1մ��5����5��ێ ������r;m)��R)8p�r;�3[�nս���N�`�  (�1&�8�m��|/�L���'?�qۙ�(,��s�H$j:<����8�U  ��6�orG��v�v��a;
�	�r98p@�ׯW��)es)��3�ݍ-��.����T__�0i������_������%]+�z�2'O�t �1��j���ڎ ��0Op/v�}hhHG���I�/mܸQ�HD����ȿ��twwk�ʕ�c  ��Y��':::�/�u�<�J=�H$�{�|(�O�3��L|dd����o��1U  ��������8���m߾�v S���:x�֭[���7����b�~�0Op�0��fxxX��Ê��jiiQ]]����ؘ���488X�m��W��;�)�Z *��~`; `�&*�G�Ɩ�^��8�```@G��4������F���|��7�����mG   �8N�1������cGG�?����b"��@4
�H$�����~���  (�\.�t:m;�u��jϞ=ڴi��( 
p��v�Z544���jN[Ԇ��>�v� �+�N+�N+����I���SUUX�.�1F�TJ)����V�}M �k��A���	˒  ��{v��J?�Q�s9���:z�h�nR07���z�G�����f���X��  �ǉJz����d2�w��ÿB�}b�o$T�D"M&�����z$��r;  (����П�w]W��?�v `<���Ç5444���Rq�~�[]m;����u��y>|XǏ���P�ߧ���ؘ���u��!�:u�J�]zc�; ��)��+�S  f R[;��˜Æ|�����Rnhٲez���|N�Pp  �t�������������H$��v
���'?��������^�K  ��z{{mG��u]�ݻW�֭��,x��#G�̹X�xڏ˅ ��FFFt��)>|X===�N~�����߯cǎ���K�ϟ��%:w �6�ӟڎ  �w�	�a��l�x.���OǏ��T[[�~�������o;  �Lc�������dr�1�^��EHJ&����ٙr]���  �L���讻�҆lG0����ѣ��.iŘ�T�Woo�������Eٽ����u��	:tHgϞ����X�D��U��j;�
��� ����2r
�sVp��U��@����顇R$�}+&�J���|  *ZL�G���7�L&�v?u���g����ٹ_��1���  ����o��6]{�c (�q�ӟ�T�TjV���\p���@���Ʈ(����Rv/��K�O����o�/�۷ێ ��������w ����>�YQn*Ȋ+���u�Y5�<oN�_   
q�������7��cS(�u&��d2�e��^2�l��  �GX�/���[�c��1 I4U>��O~������(Z	��o���ؘzzz��եÇ�̙3��y���1F�LF�ϟ����Qj�\�Ν�# � ッ=y�v @��<�=?�	�TJG��	�0k֬�=��#�qlG�����v  ��,s]���d�ˉD"��CWp��������^Io7Ƅ�7  �&���n�I7�p�� ���6����z�嗕N�~��	�6�N4*'�Ӎ�J���400�S�N����:~��Ο?�L&����\N���:}��:��G����[###��;��k�ҋ� J#�ӟڎ  (�d�#����f��
FFFt��a��@�ڸq����ʒ;w  PN:�o���������y�-7�K��Ă���0�첝  �����e�c��|�Ͷc (�H$r���lV/������:UOr��ra����b�# (2c�FFF422"Ir]W555���U<Wmm�����l6�t:���Qe2�U����65lެ��~f;
�
���O����c  
0Y�]z���g��������Q:t�r;P�6oެ��Q������U__��   ���y����W\׽����ہʡ�o&�$uvv�NCC���  ����!eg��kP�[�N��v�� �,}�}ҙLF/�����ǧ}~���   �<�S:�����u�ĉK��Ϟ=���~��i�+hc����488���n?~\TWW�Ξ=�����*�_�z���# � ï�f; �@N,6�n>�>U�+�v.���Ç+���v�ܩm۶َQV� �MƘ��������Yʡ������7��cL��Q  _
Ӷ��-�޽{C�=%P�&�D<22����gںu�ޯ��dJ����*� ��1F�LF����UUU�����GUU�b�؄7�A>�W.�S.�S6���ؘ2���٬�1����{���g�-�� S9|X���L� ���ʭ���}�?��O!<���ÇC5��t�w(�J����v����  l3�D%��d2�����[~�����L�R���������y��$��  ���^MMMz�;��ۂ���������<�k��f�Ǆy�{���v >q�,><<|���QUU��hT�H�-Ÿ�0��O�q1���/^�j�<�>������ڎ��GG�9yR�+V؎ (�����^@i��ѣJ��eH�O\��<������ٳgm�)����   .j<�L&?��O���0�Pq���?�|������yޝ��   \����#�\MM�~�a��q�Q ��t7��={V���Z�r�_��� �2�(��4��u]��{��~q��q.�a���y�ޘ�xqں�y���h�����(s�� �"}�0w ��Z��FU�/�_��rS~�ĉ�>��F�z衇����J�R����訲٬b1fm  _�J��d2��+V�}��G+jK�����S���5Ǐ?-�N�Y   �V�'�]�����v͛7�v %TU@I��ѣ:wn��
��U�"�ն# � ��i||�Ҕ�L&�L&���Q���hddD�t����,ً�v�
-ܻ�v b��a�  r'ٝ���S��w��Yuww�1 ?����#�<������  �jw?~��3�<��v�b���{2��p6�����Y   &288h;B�8���{�j��嶣 (����s���	o��h�s�� eՇ?�Hm�� *�ȡC�#  
�NR܌��.�O�L2����_�N�*s ~5�|���o���\�
Î�   ������:;;�v�b	��Jc��L&�&�9cLaM   *��s�Nmذ�v %�n�'<�����5vU�ݛfK�J�Rp��R�ڪe�{�� *�0w ��$ܥ7J�*?A�}ttTǎ+ ��b�
�޽�v�����  `2�1插��׌1����H$����aI���  0���!�JbŊ���m� P�No�(���g?��<ϻ��0Op�� �g��߯�u�l� p�S��� P��vg���������9r�9 �hǎZ�~��%3�Υ   >sOgg������E`��d�������㬶�  `:�lV�L�v��khh�}��W��Mx�LJ�t貉��$[Z��T� ���b������ ̍19r�v
 @���I�-c�r��|�믿��]� �r{��QKK��%���o;  @!�9�����>��u�DJ&��*����lg  (DOO��E�D���*�ێ�LfSp��3g��̙3�$��3R�D(?@E���k��O�c ��ÇmG   RS3��y�@���w��ʝ �����C)V��D��  �&���˅�u��8;�L~Rҟ*�� @x���َPtw�u�-Zd;�2�m�]�:�T*�w @EZ��cZ��wَ �2'Oڎ  (@�'��R)�>}�r A��ܬ��O��؎RT����#   ̄+�O;;;?e;�L�8����o%=b;  �LU�D��[�j��Ͷc (�ht������W^Q[>_�D��Rp�����W��	����`���r�QE���,4��x��rE�q9Ѩ��jE&(�9��܉v�2F���|:�N��a٬򙌼�Qy���������-ҟ~G� �a���������);6���.�Q L{{�n��}��߷�h���d����>  �lƘ_K&�k�|��lg)T 
��7�L~�q�;lg  ��Jڮ���Uw���2 ��2�]�2���64H�#S�T�A� *��jSg�^��G5��َS��U��AU����mlT�����^�pkk��q��'*�������f�O����������S�7>�����������0��

� a��.�Ց#G4~ٍz P�]�v����:Y!�y=�S*�R��  ������R���D��x�?�N$5����:���v  �٪�	�HD{��s�@0��~��Vέ��}�"$

� P�"�}�9���S�{�E�qǭ�Vռy�-X��y�T5o��,P�¯c--�͟��y�mn�㺶#��[S#����t�3�R�}|p�ү�}}���eϟW��W�CC��� �R��J�	��[�fg �亮��>��_��2���8E���K�  �1f[}}��D"�1�H��͙��D�����5IKmg  ���
)�q�jii��%ź��<��̑#rΜ)���C� B������N��?��/|�v_pkjT�d�b���Y�HՋ�QboiQ�BY=�`A`&���\�a�^6�lo�r�����)�ݭl_��Ν�عs�vw+s挼���|:�\���  vLUpw�F�=_�4e�t�̎�S ���z�}����W�b;JQ�������v  ��ZU__,�H\�H$l���o��=�\c6�= i��,   sU	�U�Vi˖-�c ��u]9�S��F�=��"�>+�r�y� �Lq PYܪ*�y�)5nۦC��{ʧӶ#��[U�Xk��/׫-z����g=yV���j��T��6����9wNcgϾY|?}Z�S��9uJ�
�ɬ�FO��� >�����*��^]-s�}RHv�PZ�֭ӦM���~�Q�l`��=0 ϟ4�    IDAT �B-jhh8�o߾k>�����3_�;::Z��쫒���  P###�#�I<׽��[�r+��)���K/�y�9_�Rq_�ǜ�*�  e���{հe��tt���߶gvG��f�R�,[v��,Q��E�8!��MM�ojR���~=�Nk��IeN��Tz��1v挼��X�̩Sj��r �&�Ko\|���p��el� PA��N�>}:��Jl  `�Yh�9��ѱ񩧞궝�j�+�'�z�uf���  *B:�V6��c���=�ܣx<n;
 ����>z�w�=xPΫ����h��� ��T�d�6�ۧ�o[G�{N�c�lGz'U�ҥ�]���{�e�Y�Ln,f;"(��~����̹so��/�އT�/�?����:e; `��y<�]�7�Lr# �V,���߯/|��<�v�Y�  �X�;��j"�X�H$|u��
���g�T�1f��,   ���mٷmۦիWێ���Op�$Ǒ��w+�o�4<\���ʁ n�o�]�v�V�/���oJ��J�3D�(�/]���v���U�t��k��s
�庪Y�D5K�H;wJ��lV߽�.y���p�d(���9Ӽg�����hj�w��S �P�-ҍ7ި�}�{���Z*��  ������~������7[�����矏����:���v  �b
����F�z뭶c ����%��Q�;�)����4��# ������r��J�߯��G���?){�|Q׉-X�x{��֮U��]�ի_�JѦ������������ڎb��ɓ�#  ������e�QR�#s���1 �Ѝ7ި��.uwwێ2+� @j�f�'��b
�/
��7�L��8�
�Y   �-���ў={TUUe;
 (Y�]���:��X��I��4ݔ7 @�4lڤ�M������4��K�я4r���Ξ�)`��؂�]��2{�ڵ�66��O _�M7Qp �Z
�f�f�\�PZ��������y��w  P������c�:�c�M�/
�������8�m�   (��!���3#�6m�
.d ��uݒ���w�NΑ#R�7��D���v ����7nT�ƍZ��c�$/�U��Ie{{�e2�g22��HM�"���SͲe���ZW�֭�#X���<O*�{o ��Mw�z࿃���m��N $-Z��۷륗^�e����5::�Z�� @�qgugg狒v��b���L&�_c̍�s   �����3��u��ێ�GJ9�]�Lc������/�t��� (��)�ޮx{��(@Yխ_�F�;������Sl��I  �p��y=���]w�p�>�2��[t�ȑ@^K��  *�M��SO��f�7�wvv���o3  @�q�����6Us!�eJ=�]�̭�ʬ��ͽ"�  ����(�j��Ve{{mG  La���+�)O��ko�Y��v
 !�F�g�9N�{���ێ   P2��<�L&�63X+�wvv��1����>  @��R)�fd���Z�n�� |�w9�̣�JQ뛍��SUe;  ��}�
� �o���icu��l�b���v
 !�|�rmܸ�v��  ��~����m-n����g��n�����  �-H�X,����v >�n�&蘅e*��tS�    �,]j;�U���
9�b���v�T_o;�������mǘ���A�   J��?��?����e?�N$����/H��{m  �r3�(�NێQ�]�v�� �R�����KZ���k���َ   �{��mG  L���{�.����\{�� B���F�v�cF(� ��pc�ط�D�/����^__��ǩ+��   6�R)y�g;FA����m�6�1 �P$R�K�Ѩ�(�e�Pp  �Vu[��V�lG  L�'��;�ʴs Le˖-jmm��`��ö#   ��1&^WW���1e=�-�b���_����k  ���w�qG�K� ����u�̚5e_��"\  �XK��V�َ  �B�Mp_�^&仧 ��qt��ێQ0
�   L�Y�o߾�+�e+��۷�Ƙw�k=   ?
ȅ�+V����v >�vf�y�|�di�R`�;  ����Ϸ�*&�������i�U����۽�v
 �²e˴v�Z�1
222b;  @YcޑL&�c��+KS�駟^���?[��   �$�Jَ0-�u5@�Y�ݡ�M�7�Y�\
�   Ӫjn��8Xɘ� �7��A�)f��^jl� ����oĎ�� @H�Igg��r,T��kc�[[[���8�R�  �7A��u�V-X��v >fk��$���jj��_4�+' e   ls"E�q�1��� ��VWO��@������i; L���Q;v�cZ�lV�\�v  �r�Hz!�H��^�¾}��$iq��  ���a��TSS�]�vَ��N˩���g�������   �s+��Y�ڎ  ��t� Lp7��*UUَ ���TWWg;ƴ�0�
  �،1������z߾}�4�<X�5   �,�Jَ0��;w�&�� ��9�]��m�I��[�0Wn�M�   
5]q�����< @�}�{K��5��N S��b���mǘw  VƘ;;;�]�5J�Rx��=���R�>  @���؎0�x<��[�ڎ  l���{���f�+�S�  &�wy��l�v
 ��inb��ws�-��؎ �ڲe�mǘw  fƘ��H$�K��%;���$Ɓ �P�s���nP,�@ X/�K27�(��؎1kLp  (\$�;�y���#  ��VUM�u�/��ʴ��N q]��S����3  @�U744|�T/^��B2����8ח�  �į���:mٲ�v ��a�W$"o��)fm��n   xS�'�K�Sp _+������y7���v ��i�&555َ1)&� ��3��L&�.�k�����k��Q��  c�����馛�l	� �����.�\���j;ƬPp  (w
� �kA-�/Z$�Ze; ̈뺺馛lǘ�  $I�D"�\�-��u6����p�}  ���=ϳ�-�y�f�1 ���蒬�ʻ��)f��;  @�(�Sp ?s���Lr̔��V���k��F��ϷcB~��  ��buuu_.������g�y��[���   A�ש�v�R$�@@���.�l�.�d��3��}  �`N��J�Qp _+���y[�̊�S �����]�vَ1���a�   |�q�[���/�k���H$����Q��  :?��q�F�1 ��
�r��ﶝbƘ�  P8'��e�\�v �
9�����C�P�֭Ӽy�l�x�QnN  ���D"Q��E;�nhh�s�q��z   A��m	���:��U���Ef�V���1f��;  ���=h9��q�  S(d�����.X �|�� 0'��hǎ�c�w  �79�SWWW�ߋ�zE9�~��Wc�[��  �~ۖ0�i��Ͷc _��2�w�N1#�  f �wy�� �)m��ٹ��� *¦M���mǸB:��1�v   �p]��~z]Q^�/����X�  P)�6�}�֭��b�c _�%��n���Ō���  
��]�ʉ	� �o�*���ˬ_o; E$�֭[mǸ��y�f��c   ��1Ʃ��y��5�c뎎���1ۊ  ����i�.q]W۶������XLf�.�)
�w  �y�ݣ� ��VUM���$3�]'��� �����UU���r�ێ�   �9���������u�|4�8���k   T"?Mp��k���`;� ���Ls�mR@��Lp  ��-��ێ  �JP&��b2�^k; UMM�6n�h;�R���   ��D>=�טӱugg�KZ0�   ��Oܯ��:� �o'�KRC��Ȃ ��    8B^p���N  �B!�}q6��k��j�) �访�z_��f�;  ��tvv>9���;>c�����   �ltt�vIҊ+�p�B�1 ��.L��qG 
PLp  @��� ��	�wו�}�� PMMMZ�z����iGg   ?1�$�1�>D��;;;;$����   ��/ܷm�f;� s|^�1�ˬZe;ƴ
��  �7�\�v�x� �V��i�gSV��m� ��ٲe���0�  `Ru���4�'Ϫ�����ǌ1�>�E  � ��؎�x<�) ���wI27�d;´()  ��fmG����.J vnUմ��}6�\{�� PZ+W�T�On����+   �����?��gu��ĉ��f�   @c|Qp߼y�\.��� |1۶���ڎ1%
�   �{�]��� �)�~�{]] v���pG�7o�C�422b;  ��Ŏ;���g�T0Ƹ����l  �t:-��f���= ��	�v찝bJ�  
gr9��r(������n6o�0�  ��/C���  05�u%�H�������%��?p�f��  ?��Z�l����m� p�(�K2�vَ0%JJ   ��w��#��ܪ�ic�l��H=���Z�r�����  ����럞�f\pw��f�  ���C�}˖-�# � �)�/Y"�|���b�;  @ἰOp�# �Z�w+gT�/�ij��2 Xq��ڎ@�  �01�̨�>������E  !�����Y��j (7s�M�#L�)�   �3!/��5l� ~V�H6
' Bf��ժ��[c��  P�ڎ��'g򄙵�]�7g�   �FGG���q�FE"� T��Lp�$s�uR,f;Ƅ��	  P8/���*
� �s~-����0�@ȸ���7Z�066fu}  ��p]�c3z|���'>q���'  !��6X]@ep'PwUW�X��1)n:  (X�'�GjkmG  L���*�qe?��n���h� T����[]��5A  � Y����@�.�7�t�.  @��<���РE�Y[@�T���m��r��  P���a���� �V�.m�>�b֭+� �����?���=�S.�7�  ��>���{2�\)��Y'  ��6��
�����l�$��؎�VLp  (��<�C^pw��~ pI���:K=�Y���+���]�����t���   ��B'}Z�Ww��.j   Ae��n{+F �#�wE�27�N�Lp  (L>���<�1�b�; ��/'��]+�e����lذ����  
�H�d!,�(���g  �L&ceݦ�&-\���� *O ����#�E��  �.74d;�UnM�v� _+t�{9Ϫx=r---�?���m�  �w�i��d�$1.  `l�7l��B* �	���a�TSc;�(�  f|p�v����mG  L�w��q���\��o���	�   3R��3ϼo�2���E  *cccV�]�n��uT�����\{��W��  P�w�  �(t�{٬_/��n� �kÆ�֦�  03�|���{̔G����/ic�  ���	����Z�pa�� ?2[�ڎp
�   �a�;w �;�Mp7kזi% �y��i���V���.  @�m��Q�Ԕ�|>�;*��i   �"�͖}�U�V�}M �-��u�⮏J宏�   ���А�VE��lG  L�O����L[�� �����|  p��y�y�LYpw�狛   (��e��L{���8���   ����n; `nUUA�+�؀+$w�K� *���ٸ.  P��Oz���Oz��%E�  �\���E"-[���k�ߙlG�����  �n���v�b�Ͷ#  �Qh��,z WX�l�b�X��+��   �-�L��싓�GFF�Ki�   T6cL��˗/W��$�"s���+s�5�#\⫋�   >6��m;�UQ
� �{~��ݬ��  �亮��P�  f�q�ߙ�k���y�4q   *[&��1��k��r |m�"i�<�)���N   ٞ����� �Wh���cZZdJ�
 ��kf�  f��}a��>��EƘ���  P�l�Ģ� ��w�G��   �l���� �i�e�6�9a ���kf���  �Rc>��3K&�ڄ����'K	  �r����u���F5s &d6l�A���/  �-�S��y�)��� ��c|
� 0���F�+�ΞLp  ��|>�щ>?a���Hi�   T�l6[�����T��i��Y�Nr'<�-+�\�  ��^��lǰ*��d; `N��KzV%�Y���+ @��\����1�  `N&쬿�*"��cV�>  @e�d2e]oٲee] ��Z��_��  �.��k;�uU���\?�ľx1� `
mmme]�	�   s�����Ǯ��[�z�p��a  �Y*w�}ɒ%e] ���`�7�  ���==�#X�����؎ ����e.n@�,-�Гr��  Pa�'N<��O^�	c�{ʓ  �2�sJC}}�ʶ�pq��n�]6~(��    ���E�lG  ���{)Ϫ
� 0���:566�m�\.W��   *��y?��&:��Y�,   ���ro� \*����n;�?Lw  𹱳gmG����  0
9�/�YǑY��T� ����r���a�	  �l9����GމD�YҼ�%  �@�܆��; ��Af�|�(�  L/s��VUSV���z�?�TSco} �r^C�<O���e[  ��߷o���8�nhh����  �<���V���~�L�  (���-� P '��1%��ti�^ *J������   @%�<�������1���  �<��PUU��e- �TI[��U����  0��ٳ�#X�� �aq��Y���� $---��be[/�˕m-  �
���s����2  �H�:��x�b�6��P�*��.�w�[�  ���)��k;�UՋێ  (��	��� ��hI�gRp  ��+:엮�c\I��  ��VkkkY��J`-��Q�1   0��s2�g;�U5� 0�����4����y�g~�_���g8�C%Q�J�(y�^�k;~�N$@�dÈ8FbA ���ȉ8�"F� ��I��țc�s���]kq��cuߢ$��x��9���]��!Q��ǐ쪧����%9�~�$�ͮ���{6�Y������������� �FY�m���?��M��������?�L �JUܯ��J�h�N'��Ү ��J!�,���#Y�}۶��-}��ڶm[ek�� pu�������ƹ���=�f�H  �2*Y�ʩ�x*���N�Hx�w��  1���֭��vS� `��q�_ʮJ�EM�6���n�; ��˲��.��~���� h�*
�N'�n�Z�: mR\�c� ����c�����o_�8��G���pe%u4(]������<m�˖ML$Y�Pp�,[�n�N�y�����; �H��|��~Kۦ� �P��[�l��D7Q kǎtk;>���WW�䣏Ɖݻ�����#�#��\}� \�Tw�.Ϲ�Qǎ+}�*� ��[��`2"�(������̧� �ULp��HE`|��!��������r �ǙW^��_�b�s��18s&u����e��#�Uɲ(��fԯ
�z۶m���n�; ��˲l�(�N�e�dD�����~6�I�  �Pńw�+0?�qcD�"af�; �������~�|��Q������ �Id������~]���Ꞛ	�  W�(��?�����F��'#"��_O�	 �5Lp���"{����Upk��c���N���Q������� �I
������; @��ÿ�
��a  ڤ���[���@Q��0���o�HPpOr���<���ś��{���������7�� ��X�u��wU6o�+��-[�T���; �hLLL�?�
�H� �U�</��;�N��ϗ�@[[�D�Y�	� c���;��o�F�z��Q���t�1}���c p���K~���6������|t:����U��#m    IDATq�3 �8(�ⶈ�
�EQ�9 ��pX�����E�$`�+��w��r���_���;�:
� 37�����I�],,T�&@t:��������R�)��  ��>"�ܕ��  #R��M&� )��,	w Jv��ߎg~�W�ہu�p�-�# p�RLpWp�r���r?  ��("":����7�{�� �zeOh�b���Dw9�ño~3^��"����Q�Qph�u<�>�{̛Yp��e�; �hdY6���~cgÆ?�: @��=�A��JQ��Vlz��33կk�;@�߽;^���2�� u�afo�5u .W���وnw��0V����� 0:6l��N�e?�: @����E+�Ql�R��&����={�_�u�v��̘��J#�U�'pU���V� , �q211qO'˲;S h���
�@U�Zp��[�_�w��Z;u*��G�(��˩� �A��q�� ��;@}lڴ��5Lp �;;��K ��
�@k(���������GS� jbn.��\�: �i=;&#�U������
�G� F�(�[;�N��A  ڢ�ͫ����� �x���ƒ{�qc���c� �s����8����c 6��O�� ���qR�HwT�	\�*�)� �N�e;:EQ] 0"����ן������R� ��6�S�^��� 4�`q1�����:�pswޙ: %�J133�W?U�_Sp ����H0� ���޼ڰaC���Q�,��ͥN @���S��:�:�p�wܑ: W`=��tGž0�U�)�a!w ����D�ǽ F��ͫ�7� >J�}4Lph�ށq�K_Jh�ک���\���H)� �ԆNDL�N �&�m�Ƃ{1;[��
� �����Q�q��	� �e���wS�\����y^�� ���NDtS�  h����&�Ukc�=�w �c���x�k_Kh��֭�ݺ5u �D��¾0�Us� �Q�:Y�# 0"eAMp��ڂ�%nD�Zf�;@k���"_[Kh��;�L���t7%�"��p��.��r/  �,�&:EQT{W ��Lpڦ���݊3��P@y�K�# -1w��# p�.� �HwS��#<8p��"�ʽt �D���:Y�.; ����y5mRP�<�SG(G�'b��h�Ճc���S� ZbV���F��R�C� -U�=6w ���Lp ������>�G���^T�~��r�v8��C�# -2w睩# p�.q�?Ҋ�=a���|��; �He�2 ��7�܁��vS~r�����w��8��#�# -�ML��Ν�c p�.q�?�q��F��{l��K HD� `��޼*{��G�u�{Vu���+�Xz��)�����'�3=�: %Qp�w �fѐ ��7�&�,dD{7�
og
� ����[�v�d�@Kl���� �
���Wp�w �fQp !܁���#����2�� ����3�# -2�kW� \w��)���; �h�� � eO� ���n�Wy"�	� ���쳩# -b�;@�]j��HwS<80&� 4K�, ��)����;P�<�̱����T��܁�ɲ�۹3u
 Jd�;@�L�<�D�
 `�:�z� ��+{���>��w�����Xٷ/u�%6�|sLnܘ: W���~��;@��� �,R   \Pk� p���%&���x�=�# p�*-�+L�D�tF F�(
w �Q*{�J��Zk��խ���μ�b�@���# p����_�N�}��^� ��Ȳ,:�-+  $Pv���P��(�Yr����� c��K/�� ��§>�: W���#��W��>@��}��w ��2� `�܁6j���n� cfI��lr2�v�J��t�	�#�	h�@
�  ��� �9ZY2j���*�޻m�ĉ�=�:�sw�����1 �Z���c�wCO FB� �Y:Y����  �FٛW��	����?S #K/��:�"��d� ���f�c�-ܗH��!R
�  #UtZ9�  �N�S������������B����^z)u�E��A��y�"�� 0Z�  ���S���k�{O�'b(�4֙�_Nh��O:u F�"��q_ ������  F�w �*{�{+K�@�q�{V����&�Pog_y%u�%fv��ޚ: #`�;@�(� 4K�, �1S�����j��p>�|�fe�����i���G����Ė�~6u F�b��#�E�'0e�cSp -w �*{�j��B&@D'���vz@#�}�5����l��=u F��	���)� #P�=6w ��Rp ��7�z�^��p>m���-/W��r$@#�}�����ޱ#>���1 ��"{%e�d����!R  ͢� 0B�N��܁Z7����ʗ���� ���믧� �Ď_����"���P(e\5� �E� `�&&&J}}�%��6��HPp7�����ٓ:���6����c 0By��þ0�U+{�T�� ƍ�; �)�mTE-*hg)&���!��P��wo�@��w�nL�Φ��eOpϜ�	p�� �E� `�܁�j�����	 h�ޡC18s&u�᦯�>n�;'u F�B܋0�����Pp hw ����,����a��������y���H2��E �b���SG Z���O�33�: �v�	�]���pU��~�{ܝ�
 �(�t 0Be�#Lq�h�ww �ᬂ;p���sq�_�K�c P���$e�dN��*����� 0Z
�  #�eYdYV������>���i�{�8Q����@}��ۗ:�`37�w���: e��>Ii�'���J��� FK� `��>�P�H�U�S��� ��Xy����������ߊ����Q (ɅNj+m�Ğ0�U9}�t�k�} `��t 0beOhPpRhS�=;y��EMph��7�Lh�lb"��w�.�v�L�2)�4�	�  ͣ� 0b&�mԖ�{����U�n���(k�NŠ��n@�t:q�o�Fl��gS'�d�Op��#K���
�  ͣ� 0beo`Uq�"�G��F�8~<ͺ-y@ `\��z+u�a��ɸ�������ϥ�@.Tp/u����+�� �<
�  #�eY��o�;�Bk&��<�f�$�p���ۗ:� ����ݸ�����Q �J��#">�b
�  �3�:  @�LN����ٳ��yt:�U�SE+�{�'������qa�;�^���?�[�n�5u *t�	�^�|pE���byy��u� F��� �*{+�sS܁$Z1�=Q�=�"ͺ \�w�R�,n��_�������0��Sp����,�	� W��{j
�  �e�; ���=�="�ĉ�y�������pSSS�c\����4+�4��}�# 5���[���Oc�O�T�( �P��^�X�T�4����+Y��{�  u�� 0bU܏;��~{�� |�`0H��>�d�]@�y���O����뮋���ߏ~�"3�`|]�!���ǎ��@+������V� ��Pp ��
� UK�U[�lq1�̙4������G�硫���wĎ���㺟����0��쏔>��{w_c�ƲWh��� 0Z
�  #V���;�B�������6��1z��� ������/�����??�c�� P'�&�GDv�X
� �E� ��� F���S�N�p8�	G�jz��s�p����c5�@��d��pCl�瞘�ԧb�g>�;"�RG���T�㽂�m�U�@;���XZZ�d-w ��Rp ����?b�yǏ��۷���9�A�jK�r"���P?
�7���+u(M656��ƍ1�eK�\w]D��: M�p�{8��;v,���f��n%�  �w ��jBñc�܁J��B�)��=�����Ŭɠ  �u�	�
� �s���Mw ��2� `Ī��Q�@DDQ1��M����G�-_4�� �q2�ܳN'fv�H ���s�_DE�'λ> �W彴�� �w ��j��;�S�: 4RG�"ّ#)�����^p����: pA�{�}��K��|�nU�K3� `�� F�����Ç#7��XS���I�7��9V�I!���nJ ���w�_�nIv�`��4�`0�#^�+� ���; ��UUp_[[3��\S�Y�{f�;@#N����r�Im����  j�?�k��(��ˑ#G*U��A �q�� 0bUn`t3�Xc���%]�w�f���&� \�yb�t����*Wh��_�� 0Z
�  #6==]�Z��l-����O��8y2iw�f��|�� p	�y�F*�-9{6bq����{h�N�w �Sp �*�UO� hb�={����o���; �%�kk���wK2f\TQ�ܕ� FO� `Ī,��={6M�*TE���1.K�o_��;W�ÇSGHn�RG  ���<����3�O .�ĉ���*[���V� ��Pp ����J׫r@D���`�����P?��GSGHjbÆ���O ��>z�?����m�'pQ�t=w ��Sp �*'�GD0��X�&��z�8��h�C c��D�IM_w]�  ���k�$W�ǏG���be�FPp h>w ��z���}�*]�Iܳ�^��+���1&�4�ژܻ
�  �4��?��$�$y��)V���(�͊�#� FO� `Ī.�/..�ɓ'+]ok*kg/��:BDD�;g�^p�Qp ���^��)���ѣGcyy��5� FO� `Ī.�G��T�Q�_y%u�����w0��<��N�N��	�  ���Sڒ]���Q�V���̦��+_ ��� F���F�S��,w�J��0u��9|8�.'\(���کSy�:FR�۷��  P��Ovf�ٳǎ�Z���Lp	�  ��� P����J�ۿ�&*͖�y#J�u�����n ��Z]�Jh�w �K��)m)wH2�O >duu5>\��
�  ��� P��7���a�߿��5��ր�v��˩#���@�>�:Br�k�M ����""�@Y�)� u��oF��t������ h;w ���԰ϴ�B�?5�ߏ�7R�x�	� �7XZJ!��͛SG  ���#�����S� ��T��Lp =w �����F���@��}�{��5*��P&�GLnڔ: @��(�'����>����(��7lؐd] �6Sp (A����ӧ��ѣ�����OpϞ}6u�Qp���Op������s  ���k�:�N�^{-u�Z8p�@,//'Y[� `�� J�j#��W_M�.0~j=�}0��R�����_ DD���b�IM�� �.���k�8�޽�:T��ڳgO��� FO� �333I�}�W�(�$k�%����c�W����^�b�;@����Iw �u��Vp"۷/u
���<���h1;;�lm ��Rp (A�I���q���$k�gP��v��ө#|La�;@�ΞM!�Ʌ��  ��C새��Fy_�pj1@�߿?�����?77�lm ��Rp (A�	�i�`��ZK���Zd/��:�ǘ�P��J�IMmޜ: @#���^�+�7ވ��S� H&���T��  �L� ���EQ$[��������S|��;@��SG  h�s������0��{S� H"��x�גf���M�> @)� � �F���R>|8�������g�I���]�ay��:BR��#  4¹���v��9�So��V�^�OMM���d�� �J� ���"|�W������{���^J��Lp����r�IM$<�
 �I�:Np��x������M`<�I�����t�� �J� ���"|��c8&� �_��z�ɞz*�����c�;@�WVRGH���  ��{���{�}8��� e�����3 (��; @	ROp��z��k�%� ��:Mq�}4u�Rp���O�̦�RG  h�|m-��r�sϥ� P��_~9�O�4� �
�  %H=�="���Ou)�g�E��T$����5�7-� ֧X[��~r<q"�C�R� �L� Pw ���ͥ����S�N���\m
�?�:�E�{i�	��0u��� �'_[�~�a�;0.�9G�MC� �$
�  %�������������
������][�x��).*7���ƽ��MM��  �����gO��j� �{�RG��z�� �F
�  %ٰaC���/F��c -6�(���g��le%i�KRp��q/�w� ֥��c0��WR� (���Z���˩cDD=Nu h#w ��ԡྼ�{��Mh����s˲GM��z
� �7��n7u �F��Q�O��sϥ� P�={���t�0� �,
�  %�ˆֳ�>�:�rIo$:�o�[��� pi���3� �e�	���١C�S ��g�I�}7nL ��� JR���[o�G�Mh���;>�l�ˡ�� y�:ARY�V1 �z��db�dO>�:@)�~��Z�����K ��ܵ  (I]
�O=�T�@�%��~�tdy+�� ��,K� )c �OS
�����N�N0rO�������  ZI� �$u*����+����:�R�� ���|��CE���{%
�A���&&RGHʿU  ��kJ�=�3 `�N�8���K�CLp (��; @I괡��y<��өc -UE��P���#�T��U�Mp�=ww �K��<����^x!�^/u��y�'�[�� ʡ� P�:�#"�{��7e��8k��G�XY�tͫ�4P�^p��[ pI�^/�A�"�}6u
��X^^��_~9u�����n��: @+)� ��n�~��?�|�@KU� M�G硇�[o�&��S��d�I)� \Z��k�5~����a� W�駟�a���6lؐ: @k)� �d�ƍ�#|�SO=y����P�ܳg��8y���F�i7����Opw� �%�z�țv�����M<�\�~?���
�  �Qp (I�KKK��/���P�ߏ�(�_�(��o��ΈyEͦ�a�>��0� ���8�=""}4�����~����z�c|��; @y� J�iӦ����G���@�E�
n�fO>q�P�딡�7�����L�I�� pqy��j�E�⋋���B� W���ǓO>�:�y�q� @[(� �dzz:���R������x���S� Zhuu���<�(w�)���ĘO].-��  Pk������G"�_O<�D-��G(� �I� �Dsss�#��c�=Vɤe`��K���=�xd�S�e2��:c^p_;u*u �Z[YY���{�g�Ff�	�0�^/�z��1.H� �<
�  %���M�Ξ=�>�l�@˔Zp���o������RG �"�}���; �ŭ��4�����"krI;�?�x�U����B�  ��� P��Np����~P�MA�y�A�y^�kg�>q�x)�]�B����� .fee%���./G|4���J�5�� Pw ��yckee%�y��1��)���� ��Oo���WWSG �":
�#  �V�������#"{���9��k �M�6��  �Z
�  %���O���XYYIh�2n8d��nd�O��u���z�# p�5~8�
��[ P��{��m(����%w�;}�t#�4-,,��  �Z
�  %��������x��S� Zd��3g�ӂ��C�jmŗ���>Q�c  �ҹ!!m9�-{≈���1 .h���1SǸ�,�j?�
 ��� JԄ��?�|;v,u�%F]p�|�k-�|n�;@�M6�{��� KK�c  �ҹ�{���8Ɉ��y��) ���ߎ�_=u�K�v�155�: @k)�*��    IDAT ��	�<���Lh�<�c0�����?�k�@+�1h��1���z�p�  �SE��{h�U��{�D�ߟ:��4����\�  ��� P��Mؔi@3�j�{��{#�b$�Um9����}�{DD�С�  j���E���D�
��y���<O�}M:ux�ƍ�#  ���; @�65h
��ݻc8����(
���OG�w�����io ��d�>��eU� �cVVV��qѲ�{��Nt^z)u
���X]]��~8u�u3� �\
�  %��������1�������SO������N*_[��W�:�05b�;@�M)�G����  j�����6�=""����6����y�G>�PQݙ� P.w ��5i��������1���_����7�q��Ճ�;@�u�mK!��ÇSG  �������ʂ��rd��~���;v�X<��3�c\�&�� �D
�  %kR����Ƿ����1��+�"�Wx�7;|8:�����C��Pk��11;�:FR�C�RG  ��~�kkk��|�Ƃ{Dd�<��|�D���o~�W54%w �r)� �laa!u����oĞ={R� n�J��E��q�p8�@5`�;@�u��6u��z��  P+��(��JQD���ݓ����C|�z��ͩ#  ���; @ɚVp������+++�c v%ܳ��l߾ч����;@�M�y�}��k'N�� P-�����ĉ�<�x���Y\\�Gy$u�+�� P���  ڮ�������w�?�3?�:
�P�~?���,����٩Sѹ���S���z�# p	�m�RGH��޽�y���1��G���[o����,/G1���LL�����B��v[Lnڔ:& 5��! E['���裑���σ@E���\Ѱ�:Pp (��; @ɚ����/��w���rK�(@E�~?������ٟ�iD���ED��?@t�oO!��{c�O�D�pU�Ǐ��k����^���_�3���o�����n���;c��xl�ɟ��O~2��0\�q������e����yd�gQ��/F�sh��z饗b�޽�c\�n�6lH ��� J�����x����_���v��� ������{�䓑��b��Rp���;RGHne߾�`݆�˱�o_�ٳ'�_=ξWj_;y�_s�ĉ8��q��G#"bra!�������\,�؏�*: ����cPp��8t(�瞋¿{@����c��ݩc\�����  ZO� �d[�lI�-..��������/��4��:
���bt�4�)����M7����rC���bE�Ç���[��o_����o����E���җ,.ơ?��8�����7�ʯĵ��\t��J_��Ξ=��_�k��ߍ��#����w���>H��#  ���; @�6o�Y�EQ��\�g�}6n��ָ���SG���GQ�]�H뢈��0�<7��h8&7��l��SGHny���8��]٤�c��?~<z��Go��Xٿ?V�|����z+�5)�,��{~�7������������o�-�?h��Np_[K�$�����w_��K�N�4@�<���gϞ�1����|�  �g� �dSSS1==�^/u�+RE<���˿��1;;�:� EQD�ߏ����~=۽;��_�8U:�2���fn�!���(���Q��8?�����tb���c��bÍ7��1�cG��xc����m�".��G1D�С����
�y���W��������Q��k�[��SG`���yO�+��i9z4�G�ⳟM�h�S�N��ݻSǸj&� �O� ����-�GD,//�7�������Ob8�����ܳÇ�s�}	���P��dt��.VL%�<�����;x0N?��Ǿ��v?^~߱#�w��뮋�5�$MJ���X=z4V��#G~�����;t(�G���ᑕ7ߌ��?��~��b��zd�#0"������������?���(n�)u��<���?�-xXH� �|
�  XXX�w�y'u���o߾x��g�ӟ�t�(@���f�`����#��%���n�I�}�~?V�|3V�|�_�t�ѽ�ژ޾=�����_w�|�1�u�BpC���/������ñz�p�}��~�PWVR�L�ȗ���Ÿ�����t��� 0+�w��k������#~�W���	} ������ÇS��͛7��  �z
�  شiS�#�{����c۶m�� ���EQ|��Η�q�P�Ti|��8��馈�K���~?zD���~O���Ԗ-1�ukt�o��֭�߻۶Ew۶�ܼ9�6o��M�"�&52E���ԩX;y2�ǏG���X;y������ɓ�v�D����'#o��Ų��x�������-n ��ٳg����6�=""Μ����ٟM�h����9���lْ: @�)� T�-���a|��_�_��_�	7�u(�"��~L�7�k��T�����Jc즼4Ԇ�nJaly�~��쫯^�{�N'&7m��͛���M�br���n���7���BLm�7���������;SS������pi)�c����/.��̙w|���S������[������o�f�������z�k��=���Wc�ƍq�̙�I���zq�}�Eޢk��  ʧ� P�6Mrx�w������Z�(@C������t����'6o��"u�$��&8@�(��S���O�\�n�C��ɍcbf&�n7&fg�397F61�7F65�������N����+,O��E��|���~?��Lw��D1���׋�ߏ�ߏa��p��rE���w��һ���./��̙��\Q�^�|�+1s�q˯�j�( \�Mo��	��yǎXݿ?���SG�(�����c�k�6��������1  ZO� �[�nMa�^z�رcG���h�(@�z�ؼys|򓟌�+(����;@3L�xc��X��G~�D��8�:
c�������㎸����Q �g.0��(��.�O���w�/��R>����<��ño߾�1Fjaa!2'6 ��s�o �j�����o;<�:� kkkq�w���|L�̤��L��a�*@�m�馏M��,E{����U�� �t�	�kkcz*]��D69�n7n����q��ػwo��?Hc�Lo ���; @�l��N�>z�y��w�#i�K���k����LO'N���w�ڛ�����Oh���3���Wph�~�k�Ҟ�������������ǎ;'��ԩSq���G���6mڔ: �XhW�
 ��&''cvv6u��[ZZ���/r7������n�)Ξ=�1���+�4��Ν�# -���3�����c pΜ9s���(�������ϯ��zO�������_�r�[�`Ж-[RG  
�  i둅o��v|�{�K����ɸ�;"˲ܻ��'~����7u �fV���������J�u:�q>���z�#�,���n��1?�8�o}�[q����1J�y���  Ƃ�; @Eڼ���O�K/��:P#�N'��Θ����w�����Y�1��9��RG `6*�#���������c �EQ��������C���˙���;�3&''$���k����[���  0� *��#[���?��?��L��s뭷���܇~��M≙��jA���܁:��#q��S� �VVV"��~}���0�������;��Q; "���?�p��Sp ��+M ���y�{DD���|���N�s�7�w���1��<���� M2s��1�aC�@���/�%���&H�ܾŅ�u��"{97n��n���0@-<x0����GQ���*˲��kR�  
�  ���~?��ދ��۶m����?��Ξ=EQ�u�=_]M�u�:������1�Y޻7޹���1 ��K��������ٲeK�ر��4@ݜ>}:���p8L�t�����vS�  
�  ٶm[��X\\�{�7���RG*�����r��>����D�a��: �4�sg�@˼����)� 5��y�.q͞��~��:��p�c1���������86��6mڔ: ��Pp �����SG�̑#G���܍{6l��o�=�,����={62�h w`�V�z+N<�P� �Ǚ3g�(��~O1����:��v�m���Pr�.��a|��_�S�N��R�-[���  06� *2==����cTf�޽�{���1�
t��عsgLLL\�{Ϟ=33��'w��ظkW�@�?�'u ���ٳ����8Op_g�=˲��'>1V��0��<��~��q����Q*�
 ��(� Th܎.|�駕ܡ�&''c�Ν155���_^^�0���x�=�MN���̩���7�L��8s��%����9�W�aÆ)E_���c�޽��TN� �:
�  Ǎ�'�|2{��1�LNN�]w�3�9�}u�˂
� �љ���wݕ:�BG�/u >`ee%��%�/��+HSO��(�G���޽���_Q��o;^y��Q�ضm[�  cC� �B�Xp������O<�D��MLL\�4�^g|/E�++�# p��GSG Z��W�Q�c ��Lo��k��
N㛚��]�v)�C�<��C��Ϧ����; @uƷU  ����#���|��R� F����w����W��W;��:�py9u .��;P�ޡC���۩c �����T������n�;w+��@���0�N�3���  ��� P�q��PE|�[��c+�-Ε�����E��b\���x�@m��Kh����SG  "�A�z�u}o���k��Lp?gff&v�����#LT����{,u��bbb"u ���� P�q.�G�[r��׿{��I����W�:Y��Z����(�;vD��kR� Z�w�@� ����GDǹ�~��7lؠ���O��ݻS�Hn��ͩ#  �w �
mݺ5:�����y�����/��\�N�w�y�U��#":c\p��g�S�Jh��	� �p9�|u��$�v5�ϙ���]�vE��A"�*�?�x|��ߍ�(RGIn˖-�#  ���nW Tlbbb$�Ц��<x��xꩧRG�abb"v�����#y���L"b0�Wk��g�ӟNh!w�􊢈�gϮ���q��>��{D��̌�;4DQ�{��x衇RG���[���  0V�DD��aP����]�N�ژ:GjEQă>�~?~�~*u����b�Ν�aÆ����{7EW"b4����W�uv=@sm��Oh�ށ�# �������|��?�����^���Ʈ]���W_����B������O��R+7n��S� �	Ûa�)������H`���+�C���?kkk���_H������뮻bf�71#"��
����P��q��'&��c���:
�"+��GED���0��.��	��������VΝ���/��R;��{�߹��{N�`��o��rD�n��H�r ��k����?�w(RG���v���y�=��W�ݣ����M[���tb�g>�:�2y��'R� kgΜ����	�#.�GDLNN�Ν;cvvv�\��p_��W��/��  Ɖ�; @�^I���|����׾�� u{���q�=�D��-���k]ĻS�ǉ�;@3m�	���ۿ?u�����kkk��{�y��D	"�-��ڵ+6o�\�������O��O���_O���Eĩ�!  Ɖ�; @�Lx��W_}5��O�ı����͛c׮]199Y����R�*����۟�܁2�H`l]���(����r�4@V��s:�N�q��}���� .�������q��Ӌٗ:  ��Qp ��+1L��:�'O�L��������o�N��K���~���I��b��Q�ӟ�6��S[������;@:�������1����ae�����o�,�J_��s�dN�8�:J��M  `�(� To5"�Qg�O��?��?����c�[n��&��y�[ry��j� \�,���ϥN���![ )���E�2��8ܳ,:�n%KU5|x�Su/�k�  �W�  i��:@��z���?��x�WRG�V�t:q�wƵ�^[ݚ�)�R���0p������O�� ������# �������=�<�}bz:�©�7o�]�v���dek�8z���k_�Z��Q����  ƍ�; @�����0���x��G�(��q�u��n�}�ݱiӦJ�����w�����|e�*� ������L�F���2�$/���������4;;��sO���V�6��`0�o|���|�}���R�   �� �4e�NEQ��?_�җbuu5uh�������cÆ���MLD�S����wMph��-[b��S� Zd������R� +�� V����q.�O|dPAU�fضm[������������_L�i��p�0 @�� Ұv��x����ǎK��믏��+����e�LO���4��w�����?�:�&y���N0V�dz{D�p��=��JY�ŭ�����'��4%�*o��v|�_�#G����DG#b)u �q�*  �1���S��_���"p�:�N�~��q�7��rނ���;0����|���# -�z�`� cei����c=��#{8)lݺ5v���n7uh��(����/~�l_�J�K  `)� ��jD8��
����7����7#���q�1fff�{�-[�����5��~�(����X��dLmݚ:�"�RG �� V��T�|uu�i�#�I�|vv6��XXXH����W���x衇�O�:�� ���ޝ��y�����e��C�p'%n")���p;���i��@�<-��E���&���i� AQ�E�E�hN�i�x��h�v9�DQ7�E�9��̜}���Ő#�8$g9������`0�9���HQ�������(�  �hI��:D��;wN����c��l߾]�=��������*Y\�}�L �K����[�e@�ԙ� ]S*��;?��	�ZO�f�:r����c����)=�䓺t�u�$��:   ��(�  ���:@�MNN�����~�ӟZG")���СC:p����h��K�r��+�o�	� k{��?S*��� !(�@��J��\���?}
��T*��{������]e}	p]:uꔾ��P(X�I���   \��  �[.ZH�f���{NO?��|���~�g~Fccc�QV�Yeҗ����Lp�x�ݵK�~�W�c H����� �	�﫺�����-��ĉڱc�u 2J��������?��� ���$g�   ���;  ������ŋz��'u���(���S��;����8�t��_.T�}&�@�����:��h0� ��T*)��|
�єN���~>|X�l�:`��ŋ�����I��%�[�   pw   ;�$M�Xd:	���ק�ǏkϞ=�Q(�˭�y
� �8�ٟՎ����c H���"�@�J�M�|�����5� JFGG��c�ixx�:
�u�fS�>�,��v�Il8  ��  `笤��ª� ЩS��������tE*��Ν;��c�i``�:Κ�ksԓ��m�7� I���L�u 	Pg�& t����T*�����3��~�\.�cǎi���J��A������?�s}���Q��#�    ��  ����)�I5;;���˿ԫ���V�e蘁�?~\?�p�6�2�������L��d��ܩ��w�c H���u H�b��0�ܜ�^oS��I����ڱc��q���ZG:�Z�����SO=��*�@�=   `$k   �q�$��TA���������h���֑��I��ڽ{�v�ޭT*eg�R���U��UR�~UkC� �c߿����u�Ο�� Ƙ� �U,7}���	��RU===:|�������lZG�"C}��z��WUw�ƛ.�`   �U��  ���f�    IDATLm��BA�������O��D�c�=�={�Ĳ�.�s4���mc
� ��\N������ 6��; tN��R���]����a����[��ĉڱc�u`�
��������c����Y   p�  l��:�K.^���ׯ��_��}����ᮞ��۷O۶m���i��U������k5� �6�ݵK���ҹ��])�� ����u H�vLo����2i'��)��h�������`Ď�yz�w���o��<�8���w   3Lp  ���.�V�z��g�����$%�D*��Ν;���'��.I����>^�v'J�Lp�����/��o$n��Lp��)
m�����^p�mxxX'N�СC����cX���q}�[��o�A����ZZ�  �&�  �:k�U�������+=zT��˿����H�����u�����ZGi�m��������<
� �H{��U�$]�/�E
�z��NhLMYG �Dj4j4m����S	)�KKC$���422���iMNN*�f& �gffF���
Cz�]�   �2^�  غ))o�Ua��ŋ�ַ��7�|�	(��|>���ڻwo����ڦպ��BPK� ��_��?��(� X�Z�W*Y� ��i���0�Zm�Vep
_e�Y�۷O'O�����u`Y�Vӫ���	��q�:   �˘�  `_��2����o���_�%;vL�T�:U�T��[o����
� �7^�װ9Z��K�t<Mw�Lp�D��ۿ�t�.���(��� �QsfF��a� �(�b�-�q�F��)��b��7�|S�җ��%�ر�:�l6u��i�:uJ�f�:>q�:   ��(�  ػ 
�P,��3�護������������5�ZM��N�>��Ԟ؂�6GC-Mq�x��
}_A��t.g �!;�74t��~�����eN4�`��i<�u H�j��V����F[�WkYÉ��F�\���W��СC���H�]�y�Ο?��'O��P�(z�:   ��(�  �;o +��y=��s:u�~�~AG��莎���:}���}��U��$���㭫J^�]Z��N� �m��A=��o���Ϛy�i�8 "�13c �]��%ɯ��v��I��(�Mn������0�����\���G��_��FGG�!ɂ ��￯7�|S�J�:V�	�   ���j   >N[��������Ok�������y>|�:��l��ٳz��ո�$����:��������x��U�l�j �a��=���i�?�'��7T�x�:��jRp��	ð�������jS��0�ŋ��G��ѣ�җ�����M� Ї~�7�x��O�#�hiy   F��   ��w%��QSSSzꩧ�w�^}�_СC����V�:s�Μ9��6H�ZpOe2J�r
V�Z�iUI#���UA�f �E[>�y}������_��j��[G1��i� ��Je�d��ry�{f�
�j���m���.]�������^۷o�b:$I����￯��{�b{||`   �u�  �$ݔ��:�orrRO=���l٢�}�sz��ǕM��h�B��ӧO�ܹs�*�'��.-m����^Q�
�G�{�i����T�~�75��˚��wT<�aN �0� �gqq����ն^/N�^p_ˍA��p�P�n�jUgϞ��ӧ�4��r�:   ��h�   DÇ���BA���N�<�'N�s����c!�&''u��i]�tIA���'������0����Y��O�=^�l `$�ӣ�����뿮�ŋ����|S�>�6��dh0� ���}������S��	/��o��jn@پ}�~�gV'N�P&��P:���ܜΜ9�.��D	t��    ���  �K�U�X�j��S�N����:q℞x�	���Y�BA�K�.�w���&�*I.�g�����%���Sp H:vLCǎ������bQ�'O�x��*�/�z���ss�t	��=
���0l�5]��N�}usssz����[o�'�Љ'400��t�� t��5�>}Zm��]��u    �Qp  �����q����ٳ:{��v�ܩ�|�3z��G��嬣���������i�3���l��$��K�]~�b 1ّm��_��_����y����/�2>���K�������\�_�*C9 6eqq����.�'�ߥ�N�.��������'z衇����ȑ#J������(�����t��Y�pZ%b�&�u   �Qp  �&A$��̌^|�E����z��G���|F;w��}_�/_��������}2�F'I��z&�Z�U�X���J%� ��k�'4��+>ߘ�^*�_���ի�ML�z�����FI�CczZ�Y� �ت��j4m�nP����q�a���A���	MLLhhhHǏ�g?�Y�������� t��u�?^�.]R֑�^iiI   �(�  D�YI���,1�ͦΝ;�s��i�Νz���u��1�%|S�%��Ӻp�>����l�޶�IRQ�^G�]�*JP��	� �M�ݵK��vi�_\�y�Z]*�_����v�j
:��
��h��Pp�M���vi�{,W�����	ð#�n�rY�N�һﾫ��ĉ:x�Y���`nnN|�A[O�D$��:    (P  DE]Ҹ�c�A�~333z饗��+�h���:v�}�Q����{�|^/^ԇ~�����<��y]y��.I%�N �\��  H�����O����w=���߸��v���Ǔ�R�O��~͹9� [a�X,v��.�3�:��knAh||\����f�ڿ��=��G�Rv���k�/^T>�����8k    ��   $�yQpO� 499���I����:p���=�GyD�\�:��z#��L�H���(]�Qp tYvdDC##z챻��O��7n�~���͛�OM)��#�r۶�w���٣�={T�qCs/�h�Ts~�: �V�T��)x~�֑��A���:B�ts������/��#G��ȑ#:x���t�r`�Ţ���u��EMNNZ�A��c    �  �䬤��:�����M�L&������:x���9-MMM��ի�|���K&�V���;)������T��t� Q��бc:����A���ܜ�7n�9;��q��ǵkל�l��eGFԷo��[n�v��ء�}����]aO�t���b"( l���bǮ8�}N:�'PZ�h6��p�.\����>>|XЁԷ��2�ǝk�W�\���u$�	%�m   �  �����}_�/_��˗%I[�l��Çu��!=��CL��j���ׯ��իW=BSJ;5},
��$�%5$�}��	� �8I��.��掠�����SSjLM�9;����Z�����j-,����0��۸"�N�gtT=۶�w�N����w�N��޽<��w�n��yJ��#�t(q|4)���x��jK�.Op���{q�S���r�=�Jiǎڿ����Ϻpܹ&|��e5�H�����   (�  D�I� ��B����{O���r��~�a<xP�����ؘu�Dh�Z�����Ą�]����Y�ahkUQ�l��7Iˊ��	� ���U���1�����rٽ��/�o}|g�9?/�R�Rz�s9�lݪ��[�UntT�[?�Sn���	�=ccJe2mϐ۶M=��j-,���q�w ؘ��Ŏ��|R��	�P333���ѩS���߯������ڳg�FGG�#�^�����nܸ��W�jnn.�k�0��u    ,��  3�nJ�c��l6WLw��rڽ{���ݫ�{�j߾}�t�\�4�jUSSS�����䤦��c3��jYG蘍��Iq�a�w ��n��u���6h6�-.�9?���rY^�$�X�W*�/��*��ˏ��E���f���hI�rJ��);<������;�2����z,34���Q�mSf`�:�$i��-���u3�`c
�BG�����Nߋ�����j5}�����%�.��JE7n��͛7u�ƍH9A���   �%�  ��(��>�ͦ&&&411!I�d2ڵk���ݫ]�vi���ڲe����6�M���innny�X,Z�ڰ��7"��"U(�"i��i���;  ���۹S��;��s� �_.˯���j
j5y���z]~�.�\V�j)�����x�T�$y��B�_z�Se��^W�Z!���m��R)e����tvxXJ����W��G�f��U$�Y�}��W*�UvhH�>e���Rf``�Ǚ�!��`��a����y� ;�JE���z��7��������p6��Ν;�w�^�رC۶m��ؘ��JeyMxzzZ���*����y�:    �Pp  �����b�����T����FGG�k�.���illL�v����a���@�RI��󚙙Q>�������|�&��m�m=6:�]�ʒ�$�ږ��|6�  �T:�4��VI����C�L�A"nV �nY\\����j��׏�ͬ�D]���<�[u]x۶mڶm��o߾�6�ʍ�q�j����5;;���9���kvvV�z�:��u    ,��  -�Y@�A���y�j������l٢��amٲE###��GFF"9ݧ^��X,�P(,�/�J*
*
��n~[�7��g3�\{����z{"l�7�  ֫��{���
���ZG�X�<O�[��tJ�x�=���wj�v"O�A���Y��ή�|&���А�lٲ�622���!j˖-F��v{�I�PP�RQ�RY^��F���&����q�   XB�   Z�=�W�VU�Vu��ͻK�R��������߯��>���-��߯��^�r9�R)��i�r9IROOϪ�f��0��qѭVK�VK�z]�ZM�z}���?��j*�J=b:.���v[v``S?����%�+����  ���	����)��-..v����j�~�e�n������rA|5�\nյ�;?��rJ��J�R���$e�Ye2IR__�Z���@�F�!i�����u��P��\^�sm��5b
�0�SI�  �
�   ��:��93�������򦮓J���f]��$o��7Yp�K�%eڒ���rY��ۭc   DF߾}J��
��:�����y�: D^�Z\\����OpO��(��c�c��f��f��b�h�v�:    >q��E   X
�4!��0)��Y�7��}}J�2��B-�W^��Q  ��t.����|�: �B�\�����L�u��b�*�X   �'(�  D�i�  �#��T*���#�7����8�I  p/��;�#�jQp�5���vI
j��<Oe6y�^�%y����i    ���  =�X ��YG��n������w  �����a�w x�V��J�ҕ�rz�{��Lp�)uIg�C   ��  ��	 �%}�T;6K����~~�6�  �$�z��X��  �����0��yn�������:*�kn ��$�|  �
�   �sN��kh��o�eڰYZ��9�^�l   rr۷[G0��=" �W�*
]{>&�'W��� ���    X��;  @��޷ </���k�fik@�  ���w�T��  �V*���V�r�=��	�I_s�n��   `%
�   �Ĥ ��?M�]����N�>L�  �[��uS�����|~���狒t�'�7� ���    X��;  @41)�����m�H��L5&�  �-�e�uS�	 ��h4T��Du�'��k�&�Z��u �Q�t�:   V��  ML�  )��m�6N�۬K�K   w�q���w ��|>������Mx�=�C% ��I�u   �D�   ��+~]M ��{;���$��v��c�;  ��z�n��`��; ���}���?���3mJEI_s�.g�   �n�  �)��� �K�4�vo�Ʃ2N�  �n��a�2�f�fSA�_ �F,,,(��?���t��I_s�.��   �n�  ��u  �� ����1:�����s��O�  �n�T�'�>S�`�0���`��~�f�Q�i�{QD��ް   ��Qp  ���� DC��L��fi\�@Lp  X]�u� �R�T��u�v���R��5�I�gI^o�.I�C   �n�  ��u�  �!�n��,�J�����Gq	  `u�>���� +��y��uyz�$�~�Y��� ��9�c9  �9�  ��#I��! �K�ɝ�,�4v'�VKA���  l���)��'�ժjFEs�Z5yިH��ǍF�:�h8e    ���  mg� ���R����\�,)�ȕۋ)�   wK����� ����.I��ܳ8u/J<ϳ�  ް   ��Qp  ���� �����$�a��  �ݒ^�{�� @���eÿ=�'���i�r9����6 ��c�    Xw  �h�;�  �%y�{��O�tg^�ơ�W*�   "'��g�TP�[G �HXXXPڝ�8\p�8p�w �nJ��  ��Qp  ���%�! �J�[*�L�
LIQ��c�;  ��:u�O\��@Ahqq�4�_���p��B�=�% ��{�   po�  �mQ�� l%}í���Q��{�G�  DU��{�hXG  s����}�4�˧��PpO�@	 k��u    �w  ��{�:  [I/��;�iZ��u�����   "�S'��EH����0��u�oJ�ZG�0�o� 	g    �F�   �NZ `+���CC�v�hOq�JQN  `#�w� `�T*Eb-įV�#�Iz����� $_қ�!   po�  ��5�  l%}�{�7M�Zڭ�"&�  �-��XG0���� �����uInOp��0�(H�Z�5��h�F  pw  ��{WK�L ���ԲN�v��H��4w  �U��޺`�; ���e�#r�����#tw �NY   ����J  ����! �I��[7��.k��5�B�:  @����Q= :/*��%�g�{b%}��59i    �G�   ޲ ���$U:�,��w  �U8>�]Ao��Ϋ�j�Fhj��p�=��)����u    ܟ��   ��c�  �$��ޭ�`%IaW�i�(�  �-�����# ��(Mo�$��[�#��	�I_k�@yI�C   ��(�  ��KZ@�AI�*Ս	��K���%�  �b��u �f��R�dcY��k5�f��Vc%�km �u    <���   �1'�u 6�>U������*_�*�#   Dw� �usss�V�U��}�Mx�=�km ��    x0�W�  b�u  6�>U����-IQ���W�
=�:  @��2���?��V��b�N8��e��2�:*�km �U�    x0
�   ��w� �H�T�nO����m�  Xs��0�N  ]���F��>�Z��`*34d�����ྚb�;  @,Pp  ��W� ���M�t��[oQᗢV�  ��J��u�|��S|����u���.OpO����N�QLp�vVR�:   ��Ub  �xy_Ҝu ݗ�M�L���S�f��
�   �$�����!�|^AXǸ��p�=;8(�R�1:*�km ��-�    X
�   ��u  ݗ�	�J����S��)�^1Ju{   {�㥳t6k �"-,,X�X�W�XG0���I{���~^�   ����  /oX �}.l�Yl�F�VN�  `���;��b~~^��[�XU�p�=��!��8+���u   �w  �xy�: ��sa�-cPp��w
�   +��(|�f�	� \����܇��#t��$ �ꊤ)�   X
�   ��w�F@���1�<�B���;  �J����O�	� ����;\pO!�6�I X�I�    X;
�   �R�t�:��r��n�y�)�-
�   +�Op�� �>�]��r�:�����u����8�U�    X;
�   ��c�  ���@�'k8̺^�w  ���R�:��L�u �|>�c�    IDAT���9<�=kt�^7y�g��Y   ��Qp  ���� �.6ݬ&�K�S�)�  �Ԛ���`*���\ �
�@�|�:�yOp�B�-Lp�4)�u   �w  ��yYR�:��i�������eŜ�;  �JM��Y
� ,��%ɯV�#�ISp�LoX   ��Pp  ������! tO��R��1:�z��r�;w  ���1���I��~� �q��.I��܇��#t��$ ��5�    X
�   ��w� tW�7ެ'�KvS�)�  �!�ZX�Na*�w 	���a�� ��0��¿CLp��#�    X
�   ���u  ݕ�{&��$���V�(%|B?  �Z5��z�uS.�'N��=���K�X�鴤���˜��Z�   ��Pp  ��$E���I�d��l�.<g�y�k5�g  ���ĄusQ�� �i~~>��%ɯT�#���){���u6 wy�:    ֏�;  @<Ŵ	�)I�,��� Ijhi�{��
�g  ���ի���FG�# @[������k������tw�9�Y   ��Qp  ���X �=I�x��t0���_*<+  @�ԙஞ�[�# @[�iz����tO�R��u��K� 	 wy�:    ֏�;  @|�b @�$}�-��)��cC�ԔT��s2�  `I��5���$H�Պ��v��{f`�:BW$}����X�   ��Qp  ���$�! tG�����������]|6  ��9^pO�rΔ�annNA�%L��{��f:Ʌu6 ��Pw�z  �&Y�    ذ���%}�:��sa�TfpP��E�������wk[��;\��*�9��ŋ�\���������k5y�ʎ�(��)�}�r;wj��!=��#G4p�RY��  iB�S}r�:����Q� �6�fS��X���̸Pp�P��Y� �=�X   �ư  o���;�&Ke#��Z�4 )Յ��T��5����UU>�H��8����97'}��򯽶�X��G�i��9��c�4x��r۶u��  ���
/�Qp�$���
�����U�f��6�	����T ��u    lw  �x{A��Z� �y.Lp�YGX��T�ԍT�N��"h65�쳚��wUz���]��R��E�/^\������)�G�j��Q>�t.׶� tF�j�x��us��ۭ# @[��ucz3���Dsa��e3Z:	   1D�   �~$�)���p.����r{�{����J~���VK����>��?Scf�k��ZX��ɓZ<yr�s�LF�,�����#��o�>�2��e ,i�̨61��Ą�׮�z����ON*�}�x�zwﶎ  m1�����W*�̸Ppo4� t���   �q�  �,鬤/X�Y.ܣ6�]�|-�E;���a�;�d�'?��o|C��	�(����UWu|\��?���tO�������C�o�j��A&��&�ժj�ML�z��j׮-���5�ժu�H�ݵ�: lZ�ZU%�%q/��7+�k3�F�p�K�   �q�  ��5QpυͷL'�KRIҐ:;��g�;��Tt��_�����u�5	Z-U/_V������߷O�w�V�����{
 ,xŢjׯ�~�[��U�~]��Y�x�E�@�����\��`ƅ�<.� ���    �8
�   ������:��r���)a�����|���b�t^������=�''��l^,4?�X��^[�P���8xpi�����}�!�?�����Q*�2��i��/�W��~]'�tD���� `S�岪1?���{vp�:Bǹ��@�tU��   �8v�   ��I5I��9 t�ӥ���Z���N�����8�}�y]������Q:�15��Ԕ�|s��S��z��Q��/�zH������ջw��==F����fS��7U�yS�����z��{?��8�� ��0��̌u�M	=O����e"�6�.�g�n    �C�   ��ޑ���A t��(o���
��u�����R*աg :��w����G
��:����U�~]��׵��w=����C|���۷����2��"h�Ԝ�Q��5gg՜�S��ծ_W��5n�t���(I��(�k�u ذ���ؗ��R�:��lDO�k'�� H�^�   �͡�  ����;�hq� ^�(�%���)��v�jɯV#�{ ���w��K_��u�X��EϜQ�̙��R�ݹsi�������Sߞ=ʎ��A��4y}rRͩ���>n��YG�:��ۧT&c 6$�%���\��`*���.��P(�9�   �
�   ����?��s\�|�Ơ�]���C�n-.RpGl�<��.��1�/՘�VczZ:uꮇ3���۳G}{������={�۽[}{��g�V�� �%h�����̨q�9=��~fF��7)�'L���� `�����y�u�Ms}���.���EI7�C   `s(�  $�O$-H��3\8>9�MԆ�&�wb�YkqQ}��u��@{�Ο�G_��� ���x~��ʥK�\����������;ջk�zw�Vn���ڥt.��� �"h4Ԙ�Vsvv�F���SS˥�f>/��uTt���� `CZ���c����8�,
�^�   �ͣ�  ���J���:��pa�-;8(�R�/r$�KJ�������l�|^��U��M7q��j����:>~ϯɍ�-���,�S�:����[\\1u�9;���)5fg�
�1A�����쬂�� �r�=��)��c��\Xc�g�   `�(�  $ǏD�H,&��2ez{����Q�˓T�4����|E��� Ї��j��XG�:4�y5�y�?��_ӳu�z�mSn����m۔۱��cc��ܩL�����E5�y���՜�WkqQ͹���Ԛ�[z|aA��[GFL<h ֭V�����|��١!�]A�H����C   `�(�  $�S���:��pe�-;<���$%JJ���u׿�M-���ut@kqQ��EU/_���e��W�o��{��Գu��[�*76���Qe��ؠ X.�7�����j��.�����z>��������TJG�X� �u�I��^�l��+w�H �{KR�:   6��;  @r\�4.�u ����[vxX��Y�h�侵���(�#�Jg�����u�k5�&&T��x�צs�����r۶)�u�r	�w�6���.��g�VeGF��+@R���V� ����o߼���Z��j-,HahXֻg�3�B �Q,U�V�c������p�Ϫ�&W�� ��d    �A�   Y^w �\����Q��,iH�{a�wDU�h����^�u	�M5gf�\�D��Ȉ��ß�������(3<����ǕJu�W�n�MyŢ�Ri�7���K�u�'�"9����  ���fcp��z�\p�:Rp����@ ���   ��  ��9I��u ��J�=N����EI��t=
k���v�u8�+��ҍ�����ae���W������Ko�=�������L����P�hȯVz��RI��)����j�U��R	�RY��Z�_��/���zܯV��뷮���;��YXXH�$l��{�%��-�es�NY�   @{Pp  H�g$5%嬃 h/W6�⶙Z�Ԑ�ۆkQpGϞ��'���<����T*�Q��O��{{�޲Y����J��O�+�J)30 e2���)�[�-y��W���ߦ��Ye��J���b�y
��{f<O��O�I���˫T�>n6ܺ�ίV�*���� X*�7��+���W*)\�� �c��;��}_sss�1:�	����	�Q�ii.	   ��;  @��$�����A ���y�}_�L�:JG�qj]Z*n�G�4���?�)�� &�[Ep��A 8a�3���  k633#���ct����7o&w �~d    퓶   ��{�: ��pa�{6���-I�6\���І� �s�O�D��q�  $^ߞ=�m�f ֤^��P(X�舠�P�jY�0�w 1Jz�:   ڇ�;  @���u  ���\'�KRQ�fg������+Wt��'�c  ����~�: ���Ԕ�0�����'��uMf�\X_uQ҄u   �w  ��yCR�:��sb�{L���6;�.�:�s��7��g  '?��u X�B��Z�f�c�r;�g����ɬ��k��^�   ����  �<��W�C h?&L�y3�"i���Z���l��K/)���X�  �[�x�: <P������Q�R�:���Аu��pa}p��Z   @{Qp  H�g� h?6��\p��EI�9���;��������c  ���А�}�: <��ܜ�����^p����Z���8�"��   h/
�   ��I�u ���ʙ�A���}�ڔT���o-,�+
�!����Rcr�:  �������fS�|�:F�yܳJe��1:.��ߨ8�5--�   AX5  H�9Ig�C h/'&L�R�?� )���e�;,5����e  �l���# �MMM)7s^Y<�\p��|-f��X[���u    �w  ����u  ���&\&�Gb�Z*�owX���UA�n  ����/ZG ��*��T*�1��+��#������rempL��S�  �0�  ���Z �^ͦ��fc^p���6v&�G�FO����/[�  �)�?��Ç�c �=A����]����Ȉu����$��&�C   ��(�  $��f�C hW6ᒰ�J�HU�	�0������u
  ���W�: �����Z��u�����|�� �i�   	E�   �BI�X� �>�l�%�X솖&��wX�}��Ο�� �s��ʯXG �{j6�����1���{B�b�^�[G �~?�   �Π�  �lO[ �>��45� )X��SpG��&��O�S  ���ؘF>�� pOSSS
�����?����u��pempHQҫ�!   ��  ��)I�u ��h4�#tE�6U}I멬SpG����T�r�:  ���4[4 ��P(�RY�d1���e�f��s?܁�yUR�:   :��S  �d�Kz�:��pe.i��Ik�5����.
Z-}�?��u  �4��/[G �U�����i�]�W�
�X�L��b�^�[G �^�Z   @�Pp  H�g� h&��W^R����U��� {�?��W  ����/��u X��̌|߷��u^�d�T�bV�������Y�   @�Pp  H��� �=(�Ǘ'��֯e�;� �<}�gf  '����P�\�: ܥZ�j��פܓ��W�� G�+i�:   :��;  @�]�t�:��se�Tvd�:BG��Tt���et��3Ϩ19i  '���߲�  w	�PSS��)�Sp;O[   @gQp  p��� l�+�p١!�Jʯ��(��む��  :~\C�>j �2??�̺�j|��tZ��]��q ��g    �E�  �?� `�\لK��(��g�#�*�
���^P��5�  8��� ���lj~~�:�)�\��`&;4�T*e�+\9p�ǒ�X�   @gQp  pÏ$�C ��6�2	>� )��㭅�nE������  pR��O;�7�c �]����{��|��ܓ��i�� ��u    tw   7x�^�`s\ڄ�I��/�~3�)���
ﾫ��1  pҞ��me�}.�x*
�Tt�X�|��K�6���$�  8��;  �;�� `s\ڄK�����{��l��݌������:  NJe������u X��}MOO[ǈ�'�gGF�#t�K�#	V��u   tw   w�@R�:��si�ǁ�ռ���o��w;
ј���k�Y�  �I;��?Rߞ=�1 `���i��o#�B�:���Аu��qix�`/��.   'Pp  pǂ���C �8�6�\8��Ҹ�Ok-,t;
q��'�`��*  @'��Y=�;�c V(��*8\��4�'�Sp/�V  �
�   ny�: ���@��Y��

�T����f>o	�W�����c  ऽ_����﷎ ˂ �͛7�cDG�+�v�\Y��(�	�I���!   ��  ��I�u ��F�K��y����E�0����U�  8�glL��տ�� +LMM9s�Z�ժ�?\Z�qe]H����C   �;(�  ��#I?�`�ͦu���8���I��Px�Z�_�Y�AB�����#  �#���ND_�ZU�Px�:����vIʎ�XG�
�@�1�  �!�  ��7� l�+q=���J���/�-,XEAU>�H��c  ��m_����+�1 `Y�����9���n�re]H�P�_Y�   @�Pp  p�_Z �qLpO�-��HRc��v�>SLo ��z��t���: �033�V�e#r�R�:���Аu��qe]H����X�   @�Pp  pϻ��Z� �1�L�riz�m-I�Eg�;�%h44���1  pJ:�Ӊo|C��ۭ� ��j��^k��[\��`�gd�:BW�a�@���:    ���;  ���� `c\�4�P*����u%IMI�|�:
b����F @W�R:����F>�Y�$ �,ݼy�:Fd�~͔����ct�+C#���u    tw   7��u  ��f\*��CGd�Jʋ�;�g��#  ��TJG~������$ ����37�o�W(XG0��	zά�����s�!   �]�  ��i� �ϥ͸�C��wjI��q�:����ŷ޲� ��i��?Ԟ�~�:	 �P�V��&���E�f�##����<�X��    �>
�   n
%1��!�6�z�d����i�j5�����^R�y�1  H����N|������i V�@7o޴�yN�:=�^�[G �q߱   ���  ��Z �~NMpwh��Ӛ��&''�u��̳�ZG   ���������g �2==�ԍ��
��d:=���ؚ���   ��  �g%��{ĔKӦ\����j6��������j�̨x����޽Gɚ����Ե���{����(�JDWHtEtEV�K$�I\�$q�Zf���4���ƃ"D.�@BPP�.CF��={�V}���>�\�սg�ww���>O�ޯ�zUwW��φ=�]������c  0�R)���������: �dkkK����1��ڲ�`ƥ��Kkj������  �1Y�    0�I���W[�{NMpw��.Iը���?k���8  �Q<^����ɗ��:
 �RZZZ���Q�#�Ѱ�a&;1a�o(���a�    ��w   �}�: ��qi3.��&덂z�j9yaaAA'BҔ?�Y�  ����.������=�� bmiiI��[�H���]��ڋKkj� Y���   ��w   �}DRU��c���qi3ΥM�Ea(�ZUnrRAhqqQgΜ�����uU���  ���N����?�cʎ�Y��;���T����^�^pg�;����$��  pw   ��%}Zҫ�� ؝v�m�o��n_{�Sp����-U�U�;��	vg�s�SĴF  �Y��9�x�+u�U�r�wS ��y�VVV�c$Jgs�:���C?�(���߭   �w   <$
�@b���S�v�_�\���Ғ�Ţr��Q"$��#�XG   ����:�������|�K�T�: ���Ғ� ���(��-��\���y�u {���&   8��;   >*�&i�:��c��;n<&=-,,����F��Q�����1  H�TJ�S�4��h���4�i�[�U�,[' �g}}]�z�:F�7��vJ*��ؘu��i6�� ��'$qD!  ��X�  @KҟJ�A�  �Υ͸�А2�����_�s�M�F��r����)�DH�ړO�[_�� @�;��ŋ��>_��-�_����u4 �g�VK����1�V��]�VʡS�\���   �w   H�E�H�6�r���J喟_]]�qr<    IDAT��Ȉ�����I���#�  0uS����T�xѩ	� ���E�u�D��kod'&�#�U���% ��%}�:   lQp  �$�����Q�  �̵͸�Ą��l�D�6��a�T*�J��}N���<��u  �"���;Ev .[YYq�b�^rz����u��rmMH�OH�C   �w   HRKҧ%��:�;sm3εib�
���n������'O�1�.
m}���1�!���׼F��E�/_V�TR֩  {�V��9ϟW��y_�����9e������Z������v��ރ.�ؚ�kkj@�=d    �(�  `�E��=��E�R��u��pm��Z���cssS###wl�n���
�M��0����O��Տ#�WsvV�+WԸrE�������vA ����#�tI�3gTܞ�^8}ZC'O*ŉ5 pK�NG�1��ܴ�`Ƶ�܁�ؐ�)�   �G�   ;>"�.i�:���P��ihh�:J_�v\������>fiiI�bQ�\��wկ|�:Bl�x����8��j��%_�t��C�S�g�e����Z|o-,P|��MN>;���yΝ�ޞ=�4�� ��DQ����RtO�(RP�Y�0��P
�@b|BR�:   �Qp  �����)��w{  [�vۙ�{nr�:��Z��H�ô� T*�t��yg������?n!�:��Ѯ���5���j��Ͻ���5?����33jLO�93���̮.> ��i�S��iN�V�̙g�?w��������h4�c$^P�)r��V�~6Sp��   �  p��w �Z���لtm��Z��+h4�����fSkkk:z�h��!���	��N|��+����s������p�_��U*�q��W�\}�93��	� \:�W��ћ
�ӧ5|�҅�uD x�FC����1�_�ZG0�w 1�&�S�!   �  p��J*K����\ڐ�:��z�N�rׂ�ԝ�722����>�B5�����1�R:�W�Ȏ�kt|\���u�;��枝�>?��������dH �q�)�ӧ�;t�:" 8-C-,,(�"�(��x�ݵ5��Ӏ�CI�u   �w   \�#��^k��!�wl��F~�*�:��ǖJ%]�tI�L�S!�jO>i!&��T<��k�s��S�oz�Z�R�m~���{kaA��$��ؘ�N����^<sF�3g4t�ҹ�uD �m,,,���X�~�b��K��u:�\t$��X   @|Pp  ��> 
�@��Tpwm�؍:���~���ZXX�ٳg0�����b��?�'�n)��k��E_�x�}Q�[Yy��~C	���2H �R����S��qN�����:qBC�|���a  񳱱�-~7�)��QΡ5��Ҁ�����!   �  p��)iY�q�  n��n[G�T>�L���эȽn��j5��eMMMP"�U����������1�,�Nw˧'NH/y�M����Z���KKj--�����Ғ���j--�S.�`%75���G�?vL��'5t�x��~�
'O*䈔N[� �X����ʊu���qx�{vxX)�Nm��$��K��C    >(�  �F��?����A ܚk�r��	g���l_YYQ�XT�X<�D���������_ٱ1�=�����ĄF_��[�z�������Zw|�����͙�F�Sثt.��Ą�G�*䈆�U��i�y�s'N(3<l �ga�T*)C�(���a�Lv|�:B_���$���    ^(�  �V~G܁�rmS.;1!-/[�0���q�Q�T*��ŋ�d2�
q�Zj/,X�0w仾�:��t>����*�>}��t��g'�_����-Ɨˊ|���w�s9e���9�};vLCǎu�[G ���ҒS'���_�ZG0������W���	�w��  �x��  �[���I筃 ��k�r�m�^k?wI�t:ZXX�ٳg{�qԸrE����iM��e�)b+75����m��KR�n�[[�:	~g����ښ�jU���qb8���NV߹͍�+�]^ڹ��a)��� H���U�q�v�sy��ck-���	�a�    �
�   ���H�)� n�ڦ\αM�k��Pd��jZ__�a&������̍�7:W�����]'�K�'�����.o}�[~/�孬toWW�)��˒�^ Qr���MN*�}�����������䧦�ʲ� 8X�fSˎ�f�/.Opwm�ŵ�4 a"I�  ��a   ��>Qpbɵ��].��w�����U�E�(�5;k��!���M�PP��Y�vBD�+����P�RQ�\VgsS~�rݭW._}?t��F:�SvlL��1e�ƔWv|���������S� 1�J��"N�90Q��ڲ�a&;>n��(������[�   @�Pp  ��<&�IIϳ�z�mʹ\p�k5E���)�Q�T*��ŋ�2iv`�WV�#��z�K�#�F��G�(�Ȯ�H�ju��ժ:ժ�jUA����[[�������s���e�o��Qe����)�o�w�~�X�� �=[XXP�ӱ�1��JEr���Z\[K��   O�n  �N��[� p=�&��vl�u�H~����Ծ���}�������J�R=��h//[G0���s�k=�.4t℆N���[-���F�[�o4���
�M����Z���A�!�VSP�)�<ͦ�fSa�s�¢�^?��� J���$e�ƔR�XTfdD��Q���ǣ�ʎ�(]((]((7>�t�ؽ�X��ٝ�9u ี�5�j5�ϯT�#�rm�ŵ�4 AI�  �x��  �;�o��/Ii�  ����)׎;Qgs�
��l6����cǎ�(��[]��`j�E/R*���cW������Z��u��ͦ"ߗ���-�7����$IQ��.�G�����A������h(
��;�����Q�l�����l̎�*���W��Ȉt�����2����(3<�T*���X�y�ƤT���LF�bQ�\N�|^�!�r9&� p ����֬c8���i��kk-���	���C    �(�  �Nf%}N�ˬ� x�k�r�M�Q��ʭ���X,jl����������������+�   ��T*)�"�(N�/��[ka�;[�   ��b'   ��� \ϵM���uS��*���(o{�0�_�(t�{F��<�   �=��H�RI��[Gq��x�=�X��y�ӑ ��K��u   �w   ���%5�C x�k�S��2Ţu3�,�A�R��0{����r|z�$�>�9�   �{����F��~��k��
J���1�ʵa@B|Lݒ;   pK�  p7[���:�g�Vp���c�Ů��M�V������>'�x���Le�Ǖ?v�:   �o�jU����1���w�X\\K�}�   o�  �,41�⦜kGg_� ��U*���?/�/�լ#�*^�`   طv����E�Nry���k,.��1�(��!   o�  �$i�:��v��(��c�����;j�}eeE5��у t|��p�u   `_� �����0���$
�n�����K�    ;   v×��! t�a�N�c��\<>{�Am�GQ���y�w Ϗ��m���(�   ��(R�T����(�_�Z�0��w v�c    �G�   ���  ����\v|�:��R�hb?�/p�{������    ���ʊ���ug��B߷�a&���k�h@�����e   �G�   �����[� ��vlj����vDA �V;��o��Z\\<����r�����    �I�RQ�\���4oc�:����u�������Y   @2Pp  �^|�: �.�6�rn�^���y��_�V���~�_#t�b�e
�   ���Z----Y�p�_�XG0��)yQ��<� �|I�  �d��  ��x��� ��Vpwm��F��%ieeE����:���Fi
�   H��5??�0��8����̵5�������H�(I   �
w   �ł��Z� @��5=�}���S�&t���4K[   ��(�����N�c�:�Op�MLXG諶�'�1��    Hv  �W� ���{nr�:��~�&��ZG06�   ��Z^^V�^���m���<�\"�l6�# �*K�}�   H
�   ثJڰ�ε�{*�Svx�:��~n���m�J%EQԷ���KYG0P  @�mllhc���8q���)�.�c�܁���$Ǐ"  �^Pp  �^�%��u�u��%){�u3��|��jZ]]������VL��O�   1�h4���l7p���spm��54 ��e    �B�   ��� ��\�>�����`�S���k���3e0���^�YG    n��<���s:V����"���
w �Fң�!   �,�  �_���u�eN��2��7�.����:�c���{ka�:   p� 477� ���:_̝wpm��;�c    �C�   ���� ���9��&���ӣ(R�Tr򂊤�
�L5gg�#    ��y�y�u�B�y
\S����x.��1ӑ�^�   H
�   دߒ�N`��±��h�Z-�F�Ah~~�Ƀ1�v��ޘ���    \gqq���b�������$-Y�   @�Pp  �~-K��u�U�f�:B����.�n�{����yEQd���z�ݯV�/�    >���T�T�c�:������ 
�X   @2Qp  ��x�u �U.Np�;�	{-�o�����i�,�us�˗�#    �V�Z]]�����~mm��	�.��1�,�#�!   �L�  p/�@҂u�E.N�rq�ص:�T�T���n�:~�:������    ǵZ-.N���i]<��54 F~W�o   �D�   �"��߭C .rqs.w萔JY�0���$����Z�Z�����#R���
w   �}_sss
��:
v�	��pq��P�;�C    ���  @/<��B%�>j6���.��*;:j�L\
�����8Je2�>l���W���2   �a���Y�>�i�"N���-S((](X��;�/ 3%�u   $w   ܫg�]��G�nι8ilG�6��0��ܜ<ϳ�ICǎYG0�om�q�u   8&�"��ϫ�n[G�x1zm�o���4����e    �F�   ��n� �k\-����`&NwI
�@sssL*����#�   ����E��u��#?f���)75e���kh��uIY�   @�Qp  @/���5��K<�S�1���icR�
�R����ܜ�0���<w����   ����U*�؇8���W�TZ��u�EI��G   �
�   腎�Z� \��]���XI�lnJQd�&�VK�RIQ���p�usտ�k��   �Z__���}�M�u3���;�    �(�  �W~C�F��\<b��{��ȯլc�R�V��Ғug_�d�^�����)   0�j������c`�:�uS����u�5_���u   $w   ��W%=jp����ԔuSq>J}ssSkkk�1�4r���ba�ӟ��   ��l69�*�:���L�84 �"����m�    �  �K��: ��Xvu�؎8�%iuuU��,�Uvb�:���Gq��  ���y������u��'�:d��Z�� �U��~�   �  �K���N�G.Npwq3�ZI،_ZZ��֖u��w�usa���?�S�   0AhnnNAXG�=��E��š.����T�  ��@�   �Ԗ�A��+\ܤ�NN*�v��l�SGQ���'�}Z��~�����OXG   � 	�Psss�<�:
z��;w ��   08�m   ࠼M�5}��&]*�Vft�:��$Lp��%���yJ }D��k�_Usv�:   @E���w���r���)�.�c�]�Ѱ� ���l   ���;   z�	I�X� \��&{��!�f�m������Yu:�(N��-����Y�   � X\\T�^���r�����vIj�Z� ���u    
�   8,d}��&]�Ⴛ����N����Y��oe��<�yJ���1ba�U��>   ܃��EU*��$]4�kYG�R\X���   ,�  p��bt�ݓ��x��477�0���t>���?�:F,��V�����  ��ZYY���u�Z���E���G��ߕ�Y�   �`��  ��Б�;�!�A��&��w�VS��X�سV����yJ�l��/��=$E�u   $L�\����u�����k��Ąu���}Jz�:   w   ��J�C ���M���u;Q$?�����J��"J�f���#�F�����_Z�   @�T*-//[��I�k�^a�;���.[�   ���  ��2+�ϬC ���hXG0�u��.��ذ��o�ZM����1���^�T���s�~�u   $����U�W.[G0��ZJ�ղ� ���   0���  �Aba8@�n��ݔݑ�M�J����%�);6��K��c���׾��/~�:   b�Ӧܐ��{!��wW�΀>Z���   L�  p�>��$w ��M�����;�ؔ�����ښu��4��[G���w��:  @|E��JE�R���� �V�N�W�fS����0���Enb�:�	WO?��%��!   0���   0�BI����A�A�l6�#��ML(�N+
C�(&:���zbuuU�tZSSS�Q��K_��}�:FlT{L�<�C����Q   ����_��jO=���O�1=�������[>>=4��'T8sFc/x�F��|M���ʎ��9��j�ۚ��S��kK���Zz�\������'��_�  ��E�   ��%����u`�8;�*�RnrR^�l��� ������N�599ie`L~�*��+�<�(�1����|�K�Js�!  |��5._V�T{�)՟zJ�RI�Ä��VsfF͙m<��$)��j�4����}��*����=���쬂 ���>����)�.�c�����JZ�  ��E�   m]�H�Q� ��i�Z�̸\p�ئ���$Qr�L��ɗ�D�G�������'?�c��}�Q   z&���x�iշ���˗ո|Y~�v _/�}m~�K��җ4������_�ӯy�ƾ���$��433#������\]C���R��kg@��:    w   �ïIz���u`�A�N��\.g��o�Z�]�����N�5>>ne z��(���7�I���[��~�w_����U<{V�L�:  �텡��W��7�~Z��]���=Me�i$���>��O}J�^�2������^`�e�:��fgg)�;��ܴ�`��5&��˒��:   w   �×%=*�[�� ���l:Yp�:d�Lgc�[dI�5CQia�{�1%�{w�;�SO��-�1b%
C5��Ԝ����Ϯ~>�ͪx/]�ȥKy��4r�}*�:5P�� �d�U5�\Q��5�\Q�'T���S�	�?��Gѱ��^]�������r{�ӱ��>�<O~�n�L~j�:��F�aT�a    ���;   ���E��f��d!8Υ��v:
�ueFG����N�=�Jill�:N��:��K�Ըr�:J�E���v�l��g�ǻS�/]��s�������}�)˿M  ��rY�+WԜ���.2=���������'���Oh���s��&��o�Nt��577'����7�'��Evb�:��V�/�,�}�!   0�(�  �_> �%��W�Z�;<�]�n���.uK�RIgΜ�� ���i�;����=�UU{L�����CǏ�xႆ/^�ȥKW�w�T	  p{���n���g�}�rE~�j�@t�e��O��μ�u��?�T&cI��fgg�n����H�񂻫�W<�S�1�A�I\=  �G�   ��;��笃 ��Ղ����;:岊g�Z�8Qi~~���=:��߭��1L�����jo�+    IDAT//k�_���ى	_�x�[��N��R)��  �/�P�RI����+W�|�5��4���/�4����~����+��L�h'���Pnw\bOG�WO�su�8`���Y�   �(�  ���*�g$孃 ��գ���ܽߜߙ�~��Y[�I���@�s�Ԝ�����RQ�+_Q�+_���b�;���/^����tI�3g�ʲ, @����Z���McoNO�1=��������뫯�����լ\�!��!��{nj�:�	
�������   p;i   �%I��j� ��pu�.�������u������(�߃c�x�f��N�N�M՞xB�'����lVųg�+�o�Ӆ�QZ   IA���5E�����O?�V��(��%��׾�����Z/���Pfd��_{����E�ޠ_$~7C�����f��Z   �;(�  ����(�=��f]fdD��!�N�se�\�����ٳgU,��$����
�1�����u���R:vL�s�T<{V��g�E�s�T8sF�<��  ���5?�����o33�����jO<����O���v�����5w��^��\�H��R)e�NQ��.@�=)�O�C   ��  �o%�I�f� � py�>75�`q�:�	�J7Ahvv�I��P<^��{�jO>i�Ej//�����G�������/^��}��p��շ��� �-x���)���j�Jj�Jj\��������Qy�1}��o�s��kQnǭ���F��q�r9�&�> ��ۭ   �-�  `�m��k.o�妦�r�����ajnnNgΜ��Ȉu�D9�=�C�}��ժ��?���_G:��M|߹:uJiG-  ���KK���|�vnN�����z�uBl[��'4��:��;ԏr;n���a�Lnj�:�� =U���   pw   X���7K:cH:��[�>l���X�]�U���)��ѱW�B�>�(��� ��Zj-,h�_���tZ��'������N)�ey o��U*�97�l�}������ӱ��]z�WU���*�?����@333j��=n$[�騳�e�L��!�f��u`��[�Q  ����  �_һ$��8�x.�so҆���VSft�:J_�Lr?}����Ƭ�$B��QM}�wj����:
���Z��Z��6>����Je2*�:��ٳ:sF�ӧ5t���۬c�c  v������ו�WV�(���=O_��_�7��o*�N��y}����,�v�Rgc���!9����f���   @_Qp  ���J�YI�����-�<�]�Nq/:X>��H�R����|��)�㖢 PsnN͹�[ޟ���Zv/�:����ݷS�4t�ҹ\� �*h6�^\�z������E5K%���uD�I��_��G?��zUO��r;���Ю��p 
�@����y�   pw   Xٔ�AI��u �\>n��MZI���U<w�:������S�4>>n'�&_�RN�Tkq�:
ƯT�U�h�o����R��G�^-�_[|:qBCǎ)�e� \�ZW���ś�읍눈��w�SǾ�������t:�����y=J�A�Y_��`*?5e���C!��5�    p�L   ���%��zw.5���Q�|̶$u�BE�E�&&&���Z*�։�AM���Q0@�0T{yY��eU{�����9��ɓ����:qB���ɓ��� ؗ��P{iI�[Naw}B2��[]��C���^���܎�r��S�Ⴛ�C!�zDң�!   �&
�   ��w��L�wY���iT.O!�(�Kݒ���TrJ�wv�~@3�|�� ��W����y++�>��-����Zx/�<�����	��Ç�T����=a�}��%oeE������r����"�V���S��t�5��׉/��inn�r;v����y�O�sy�衷Z   ��(�  ��w`�\���Q:�W�h��s����Nr�����[��Gu��/�ڧ?m�ʯTT�TT{��[ޟ��?rD�c�4t���G�>[~�~?��R�L��@rD����G�׽��n�}eE���p������|FG��?�۟�<������J�A�|�����\^3zdF҇�C   �]�  `���Nr�u �\?n9?5��Ғuܯ����05��d�;9��?J��v:j-.��}R�-��:rDCǏ+w��
Ǐ+������S�������>�Uykkݷ�իﷶ'�����)���uT��?��=�[��fggp*�������Q�r9�f��ܳwH�I   ���  �8x��_�$Q��VEJ�R�QL�.��>��V�����=j%��_�B�������_[Gz'�^YQ{e�K���=ڝ�};t����G��Sp ���ݾ����)�_Sbo//+�׭�����cj�̨x��]�h44??O�{�r�=���܁{R���Y�   ��(�   �%�?H:iH�(��j�T,���py����!E��������� t��	�(�t浯����k����*��*�����𰆎Snj�[|?|���#G�o�+;1ѧ� F���Pgc�[T__W{eE��uy��j����]^=�:-�7���.��O��1�ZM�RI!�`��NG���^3�(���=���C   �m�  ��ߒ��� I�r����ڰ�QgkK��q�(�����0u��IgO7���/�
gΨ5?o����PczZ����c����9��ؘ���W'�g�Ʈ��WvlLyN� R�n˯V�NY�����W��?�VW���P��i�&+��.���R:}���ժEQ��ax������P ��;p<I��:   @�   q��J�I��A��i6�:t�u�Ç�#����)��F�RQ:}��ҷ)�8)����=���X'ϯV�W��zl�PP��!�V��!�&'�S�VnrR��I�''���辍�+1`!h6�)�孯���)sS�5�������:�:�ln*�}��@�WV��裚��o�龍�---� �66�#�rz(@��D`�~_Ҭu   ��;   �bC��J�	� @Ҹ<�*�h��W.�x�u�ت�j���י3g(�_��+_��w�[^�lpF�j���������d��)���+;1�����s;����n9~|\�B��&@�Ea�`kK�JE~�����(7����!E8�����M���u���% ����w��ʀ{Ib*   b��;   ��%���r�A�$i4�̸>�������u����ܹs�d2�qb!](��k_�g��6�( n#
y��ϧ��n*�gGG��ގ�<{;>~���ϧ���o�M��
�[[���Bzp�b��ǝJE�֖��-�� �h�/�BA����$ieeE���Ʃ0ڎ�;r����Zp�>#���!    ��;   �eF��$��:�$�V�:�����;�o��V����̌Ξ=�\�k�$��?�������ܴ����v[���9�6��>[�S��b��%��Ȉr��J���
ݒ�А҅�������=��!�fSa�y]1=h44��k5������f�[X�yL���^�_�)l6��8&h6�����x�������葎���\pg�;�o��u    `w   ��/I�AI)� @R��u�f���J��Ζ���{�v��$�|>o�\fxX�_�ZM?��u 1��:��=��%32�-��ʎ�t�����+��w�
J=�~>��ؘ$]�X��������J�rR:���H��+�e��&a(�V����������n����z����uEA����NSo6v:
[-����^�ZV�)�+�,�� n������ߨ-Na@�^p�;<�	���|Uҧ�C    ;X�  @�|I�Ò��:�NO�J����Rki�:�	&��M������Ξ=�"��u�~H����J�:
�����t��2e�-�g2Je��KR��N_}|�PP�6=��������rJ��=�)�� �)�_�qp��W�;v:
�)�G���R�	%]���u���Ջ��^�~͜���+	��Z��f    �w   �ѯ��;�k�O�ʹ\p�ذ��8AhvvV�O����4`We��u�u��3o�u �(�W��t� o��5I^h�_����n�H .Op�NMYG0��i��>�$��u   �Z�?   軏Jz�:���>r�+��(���8aj~~^����Q̝�������1   ࠎ�I��Ǜ���a���;��5y��Lp���%��!   �kQp  @\�� @R��i�?|�:��(ԩT�c$REZ\\��ʊuS�|^�~�ǭc   �1mI���IW{�)y��F�0h<���Kn��H� ���n�   �
�   ��ߖ4kH׏]�9>����n!���׵�����I�ǿ��5|�u   8�)iMRp�Q����G<�_+g>�N����oJ�Z�    nD�   q�Kz�u 	\���z���M�^�T*���S��QL�2]x��c   �5u���͛�;z����C���Ppv�.�-�!   �[��  �8{P�}O w���]��M[o�o��P��533#�����8��k�[��:   XE��]Ӝ�U�T�G8��Lpw{�؃��=   �w   �YK��1��/�;�i�K�VK333�<�:���~�g��f�c   `�D��%Uw���/~� ���/�>l���ke�.y�~�:   p;�  w�&i�:g�z�:�������u3�o����y���vr3|��%�����  �JZ���YʕG=�4p����>���2`�>$i�:   p;�  w��k��f��(��c�I��w���6���@333�Vw;crp����P��Q�    ��I�=���ܜZ���.�8\p�
���1L�x�:�G���  ����  �$�e�}?pF��<�:���Ó�\޴?HQ�T*iuu�:J_e��u����   H������>�<S�qO�H^�l����%���˹��>.�k�!   �;��  �$X���u �\߸�;�y���
[-�kmmM�RIaZG�c�x�&�雬c    ���$���_�b���E�֖B��>�n���d�.0�   �G�   I�K���Q`���q�?|�:�)�)��Z�jvvVA�ȏ�TJ����)��Z'  @�T$�K���C33j//� \䭭YG0�?r�:�)��������	.�s�!   ����  ���;Il�+��o޺�y��fS�����8|�N��Y�   @BD�۫=|�ʣ������/�9>��52`~�:    ��  �$?�{�f�i���޼���4==�Z�f�/ο�*�=k   1HZ���J�&w�����FB���/J��   �nPp  @�|E�'�C q������:�o��S���W�\��r�2Ţ�ޛޤT��#   �ZGҊ��<w��y����t�/w��;ׇ@ w�    ��%   ����=��5\߼s}:��+�"-//kqqQQ4�?��_�"�����  �j�[n��k0���w��H\���>f   �-
�   H�/J��u n\߼K
ʎ�X�0��潕��M���+C�(��ߨ�s�1   #[��$�o�
���/O�����Na��52���  �D��  �$��b�;p6卵������j5=��3j���QL�P��{ӛ�4�H   ��$�%m�?3���V��2����s��J�r�1L�~�!p+��C    {��$   ��Ie�6嵐�G�#��ln*
���<O333��ڲ�r`�_�B�}��c   �P iUR��_4����c���H�����j�1����G����R@R��  ����  ��z�u  Nؼs{���P�r�:�ӂ ����VVV����ox��x�:   �%-o��[��;����rG�XG0��&�%=d   �+
�   H��H��u .ؼ��o�z��� i}}]sss
��:Jϥ2=��~I��I�(   裺��ۭΌ�=�^�b�:��6r|mD���u n�,i��   0�(�   �~�: l�Qp�8>�.Nj������y�u���;����Je2�Q   p�"I�����m���&@�x��6�:d�C ��\��>�   �~Pp  @�}L�Tb�N��[G0��xi�ۚ��V�^���s���mzο���1   p�u��׬�l�<��v����9�/��4��Á{�1�   	E�   I��� q���]�RGAhnnN�r�:J��+u��~�:   @[���m\T\�,��#)\/�9~���Ӓ�e   �/
�   H��H��u��wRvlL�|�:��7��*�"-//kaaAa8X�.���s��_Z�   @�՝�X������׿n	����Lp���u .��$�:   �_�  0���Z-E�O�K�����Na��M���T*���V��9�����_�ox��JYG  �=�$mH*o�G�����p���t>���us�IҌ�w[�    �w   �?���u�R�j�Z�1��>��[_�\��!���fffT�V������/��_���(   �_Ҳ��u���|���wQ�N�l��L��.>w`ۛ%u�C    ���;   �/X �����������ڲ����@�RI���u���.=�ۿ���﷎  �=h�[nOB������u�XgsSQX�0�s�T�k�>芘�  �@�   ��c��h����wx��$uVW�#`�6775==�N'	U��y�s���ާ3���Ki��   �,�T��&)4βU���<�_9|���v��0L�w5�@�Y���   ���   $Lq�Ӛͦus.Op�����I�j���3Ϩ^�[G�t>��?�S��~P�^�2�8   ��@Ҫ��u�}�Pp��^pg�;� I�%��:   ��  0H>.���a�T�ݯ��w�7�(���jee�:JO_��ox�[�>��o��8   �֖��}�D�'�T�k_�F{�^W���K�I�(��  `@Pp  �������<H������O����s�G�"=<Z���UQ�.�D(R'T�
��ǔd���� q�;��f3�8)(pT�NcS(R�yĳ���Ν����}��>�䏞陹w�ޙ{g���������<��w���s�?�&��7��upp�����}�Q���>������}���Z��oQ�T2	   �ZLn�My
a���˦c`Dy���F%ggMG0��;"�MI�b:   pU(�  `����ϛ��"����V̊�[ݨO�w�mkmmm"OV)��z�����������~�r�=g:  @$�*��B�Y�B�K_2#ʉ�I�)
��~����  0A�    ��G%}�t঱�'�	%�e�ժ�(F0�}�y����u���kv�	V*��~P���$�=8P��W�~�55_yE�k�E��/  �u�I�J��}�Z/�,�������E�=q̲���1�8�? �^��  0a(�  `���?��u�� 7�E����ld���E�	�����d۶n߾�Dbrߤfg5�u_���;�����Q��W�~�U�^}U�oȫ��  ?�����&cj�I}ۖ��ʿ���(!���c��(�K&M�0���������  ����R   D�'4(���DdPpH��J_���F��/�Z�7�سm[+++�}��
���87&����Ғ���_��o6�YYQ���~�5uVW�Y^V��  �&_ҁ��'U�O���;N�� 0Ø�$�G�eI�e:   p�(�  `R�{I�����
�Q_����Sp� ��kssS333ZXXP,�����J�{�J�{���WwcC��^�����ʊگ��   $�+��A�}����e雿�t������F���LG	LpGD}RLo  ���  �I�II�d��
�Q/w������n:�X�ZU��ѝ;w�J�L�	�DB�^P�N���﫳�*{yY��^S����Y[��4G  0�BI�4�H    IDATI-�AnH{yY�m+�ϛ����홎`T�O�?±1D�$���   �u��  �I�ǒ~G�_6�	L�HG|jY/����q���iiiI�R�t�����Wj~^���x����,�+_�����ʊ:��r&  x�X"��[�28�������j�w~��s��$�Fj��ʩ�|�6�R1�������;"�M    �w   L��􍒒�� ׍E��d��nķe�t��kkkK�v[KKK�,6)��x6��߭��}��~�%��=uVVd����++r��%  Qu�Ȟ�sG�Ýjro}��;�8��*�ے꒢�WM��_����������qLG n��ux   &w   L��H���K�A��F�} E��t܀F�!�qt��me2�q�V�XT��P��8u�W�����Y]UguU^�f()  ��\N��S���%��W��畽sG��ɋ��w�}�Y���I�����/����E|�;��v�m:pSBI�4   �N�  ���W$�M��mۦ#��x6�D.�~D�=
����������Y���)���41���*�ר�5_s��~�9,�w��e���������� �sS �y�ҰȞ{���4��S��-�)_��>�����EYǕ[�ʹ_�۷MG�p�>�}~�t����1D��J���   �u��  �(ؐ�����t�:��+��L&MG1.97��Ɔ�Fx��B�S��"!CU*ٶ�۷o+�J��4���J�}�J�}��ϓ��'{yY�������Uu���w��� ��K$�^\T�ΝA�����{W�;w��s�ʿ_�T*j��B���GZ��B�
z=�[-�1��g2���c�
@ҏ�   \7
�   ��OI����� �u�v��%�ԍh�]a�^�2����v�Z[[�����8�c%��E�~px�mo���������KowW
C�� �E�,K�%e�yF�g�U��g�}�[�{�Y�������8��߿�^���K/Ezת�گ���}�t�V*�~m�ZX0adt�w��I��!   ��F�   Qq_�/H��� �ɶm�J%�1�K�͙�`���O�=�|�������nݺ�x<n:R��,����_{���;[[�޻'gkK�֖��  DW�T���Nc�ܹ��s�)������ժ���xc��y�j����\����k
�P�X�t��홎`T:��@�x�'�uM� ��+�GL�    nw   D�ߖ�m�fM�[1D}zY/��Q�j���tt��-�E�qp��KR��TwsS��uu���ln'��L$ ��ųYe��N`ϼ�-�>��r�>���(�y��߿�D��������m�Y_W���LG�A�J�t���%1���K��4   �	�  %MI�Pҏ�\��>����7����{��ijjJKKK�,�t$\B�TR�]�R�]�z�1�Z�s��`���k��=�ժ��  ��XL��ye���Hvt�޽��̌��h4���+���|����*fY
������֫�Rp�87�����#��> ��   "��;   ��'%}����� ׁż�T�w{_�ǱF��N��۷o+�˙��+���QrfFů��\W������A�}kK��uVV���QxNA �qb�RJ��K�J��=�x6k:�S�}_���j�Z�|^�XT����YY��d����+Z��o0���,��@�pL�ӒvM�    n
w   DMO�/�gM��yQ_܍��:��y�666433���9��O0+��������~_���CSߝ���ܿ/�� �Q1AS�/��ji{{�ܩ�*��=�%�o������MG�!Q?�;��@���!&ܾ�   @dPp  @}Z�Hz�� �Uc1o�J��,��5���A�
�Pj�Z�u���#(�H(��3�>��x��l���Vo{[���������Y  .#��>T\O}|���T�t����vww�h4.�y���j���o_S���;�:++ʿ���(0īTLG0*57g:�H`�&�ߓ�6   �I�  E���-�L��y�Rss�-��m[~��8%f<�u]����\.kqq�i�J�J*�J*��ҙ����JE���`�������ˍx� pZ�TRjnN���S��SssJ��+s�����9�ͦvvv.<�����ަD.�>':�����#ʷ�H�H���?�11L�5I?c:   p�(�   ����?���A���bޱ���1�q���}�Y�10����:���qaV:=,'������m[����)��﫷���ޞz�����ȭT>Aq 0�,K��y�o�R��me���^ZRjiI�����L�tʑ��������S��,��.տ��+L6�گ���o�&�1`���g:�Q��Y�F�b���$�t   �Qp  @�����[c�01X�;�-�{{{��HLs�U���ʿ����S�@�����m�������}9��rwvԫT� ��� ��,K��Ye�����WfqqP^��W���ܜb��c�i��?����Pp��y�M�a�;DN/�;	���MG}��zYү�   �@�   Q��H�}I_o:pUX�;���"��E~\\�^�mۺu�����8�T�����c�m�7�r����ߗ[���ڒ{�vog�I� ���2w�(57�����v��vzqQ�KG��*��?����\��g�NG�榲oy��(�aQ���c'qLꓒB�!    8J	  ���!IQ��0X�;�)f����#��icc�i�0.Q*�P*���w��x��r+�vw��j��jU��=y��p �ZU�4x �,%�����UzaaXX?*���攜�Sjv����j5���_����Rss�ܾ-���+������?��AQ?����1v5�����3   0��;   ��O4���#�� W�żcQ_��E|����4���%
�q����q��^\|��@����rXzw��O���]�k5�w3���,��'>N��S\q��jgg�ZOF.����%��xCs����aQ����Ob�&L 飦C    &Qp   ���W$�M��y�R���YVd'�2�O��<mnn�P(hiiI�d�t$��,kP�������G>իՆ�w��@n�"�RL�?8�W��S�K������Ai}zz0Y}zZ�����rY��Y%gg�ω����
�p8�=����w�S����~�q`���0 �ܓss�#���a����?6   0��;    mK�I7xZ��(C�b1�Q��%�J��r�U�Q�p+)%�_�j��Z]]��ܜ����w�D�{�[�ܣ��W��_��wp�~�.��c
�@4%����%�SSJ����J����GL�N�����z��~���]�����q�U������+R�0�'w�)�Qp��H���   �i�  ����I�L�F�v���r������\d���k4�,�MG��}_���j4�u�2���H�Q�r���?��a8(�?�_���j��l*��"$���s9%���8,�/SSJ���"�Q�=Y.+��������U��� �|^�瞓��r��w�o�A�=B�z]�癎aL"���͚�12:����U�I��C    �Qp   lI?���c`�ٶM��Pj~^��6���>w\	�q������i���˲,ӑ���]����I�fspi��5�[-y������u��~���u���G̲/�,��׉b����ǉbQ���aQ=Y.�J�L�ǘj����ّg�l[x�;(�K���5��_k:n�[���`'s�P�㘎\�=I?n:   0
(�   �~N�#�]�� Oömͳ�)������r/�h:&D��V�j��Z\\T�P0	�8V*��ܜRss����qN�O���}�VK~�#���]�ݮ|&^b�X�⹜⹜���٬���`��ai=Q*)yXZO�J����|��q]W;;;�m�h��;ߩ���=�FAgy�t� wo�t��~��$۶����U�1I-�!   �Q@�   8H����5xl�|,��^w�tL �u����B����%%�Iӑ H�2�3iaቿƃ��~�5�}���q�s\��v���o6�?�۽�.��)�H(Q,�J&ee�ǥ�lV�BA�BaXZ��r���y%�yY٬���9��b��	x�0U�մ��� L�Qᥗd%
�}�Q��nn*�<�x�	�����1��L�d\�?����C    ���;   p��I���?o6��X�;���bo/���p���VWW5??���i�q \�D�(�W�������W�ݖ�`�q�8
\W���w����}_�mKa(��|�VKaʷm��?�\�S��)��z�|�Q��Gz��J��d�3Y���D� Y��nK�%��g���s9�D9=~XN?�/�HJ�鴬TjP@O$�(N}O J:��vvv���LG��i�^xA�7�0Ũ�����T�LG���I�O��Ϥb�&��5�   @�  �����/Jbl ��z�2_�u+�0�|���Ύ������LG0B���ҍ�0��xI�������Q�~xG8(�? �<��D�=���g��R�?��dΝ:|4%]:<AR,W<��pF O��}U*U�U�Q�Tx�;#_p�${y��{DD�=/�c{�����6   %�  ���I�%�æ� O�E�c��Y�,Ka��GQ�f���8����555���%r`N̲*֟]��	�P�ZM�JE�s��K/��0:++�#���ߵ,��`:���X�\ �c�C    ��2    Q���G`��w,fYJ�Κ�a�{p�p�8�<�FC������W���   <�N����U���t�]��o{�bKܣ!�#���M�����!�ܯI��L�    FG�   ��ݗ���<	�NKFx��0ԏ��?n^�T*Z]]�  0�����߿���u�z=�q.��d�}�Y�1�s����x�y�ݭM����L�t���n3�c˖�I�!   �QD�   8ߏKZ7�,
�����MG0ʉ���0���iccC����<�t  �	�P�jU���j4��\ZᥗLG0/���0�׬�������=`��O��   �"
�   ��z�~�t�(���^\4�(w�tD\����ʊ���Dx�"  }G�[vww��uK᫾�t�����4�,��u��#�
�S�����   ����   <گH�C�!��`Q�T�'�G}��!U*����u<  9��w�q]�t���g��$ɡ�>�܈Op��~�31�~H�c:   0�(�   �����st"���iQ����옎 �����Mmll�qX�  f�����=���L�NX�RI��%�1��nl���k��`��8�1�G�~�t   `�Qp   ����[�C �ԪӢ��ۣ��d۶VWW���%��L�  ���ժ���upp�0MG�R���*��s��&���E��n2��=��;�L �L�    Fw   �b>*��0��z��%r9�1�q��$�Q�fS+++���S�Y
  �~�v[+++��ݕ����\����f:�q���abE��7�'�?�a3�*鋦C    ���;   p1�%����E��}��k:�HIEx���8�M�1�sA���-//�^�3i  \�n����umnnN����[�j:�H�nn���k�5��tcb�R���c�۶MG .�%��C    。;   pq?.���E��wZjq�t���]������������;Q  �+�y����"�#s���T�t�(�O����M��K���##Cu�]�1����%�   �
�   ��9�~�t�"�Rܸ��o�݋��?Ƌ�8Z__��Ɔz���8  `LA���}������b��ܳϚ�a�s��*��q��K�Y�Q�c �.��   �
�   �����k:�8�OKQp7�4۶��������}�q  ���P�jUo���*�JdK���7�8w�����?ۨ�x�b�|T�!:    . a:    0��O�Kb�o��v�m:�Ha�;w��0U���h4T.�577�x<n:  Q�fS���r]�t��/��}�!���Ja(�b�������LG0*��8Đ��ߗ�/M�    �	�  ��{E�?5x�N�D|�;�]�I�{{{���
  �f۶VVV���E��P�LG0����5�c�D�=nj~�t���w�W��   �
�   �����aha�OK��*��n��19� �����|�MPt  �l����666���L�)��%ųY�1���옎�k���Lp?�c`?���    �@�   x2uI�t�<�v�t���,�fgM�0����j��\����������u�ah:  �A�nW��ؐ�8�㌤X,��3Ϙ�a\oo�t\1��T?�f
8ށѶ#�S�C    ㈂;   ��~V�M� �B��a��E��br!&��y�����ꪚͦ�8  �������-���ɶm�qF^��]������I�E��4Q,�bw�S�}��	I��   <
�   ��%����A�����T�'��L.���z��  �`������Z^^椶K��.�"^��DQ�3M�ϛ�0rx��EI��t   `\%L    ��J�MI68�Ž�E}���wD@����Ɔ�٬���T(LG  O�u]��h(C�q�N��{��Гȉ���Q?y�,È�%}�Cr    <
�   �����o�T28����R�r�wDI����榲٬�����MG  �ຮ*����&����wɭVMG��E���4����m������/�   �3�t    `lK�	�!��X�{X���^@4Mt_[[��E  ƀ뺺��VVV��~Ţ�h����
��t\��O������^#�@��4   w�  ���^68���E}8�% D��D���5�M�q  �(�_��3Ϙ�`T���o��o������Pp��[��   <
�   ��$}��5`\�ݦ� +����¾m�g�������E� �A���en�2��~�a:���n������#��<`�|QҧM�    &w   ���;I�a: IA�q�1FNfq�t��������j�L�  r�~///Sl�f��Y����u�pE���6��w��1B|I�'�6   ���   \��T3�آ�,��o��2 �n��{��iyyY�jUA�F,  \�N����MvS�Aɹ9��c����{�������1R|�W��38�iI_0   ��  ���'��H�ϒ��w'�e �<��jwwW�����ߧ� �k��Z[[���:�SnX���\&�O��ܣ~��Yl�f��I�0   �$	�   �	��J�vI�3����,-��`��2 �8�~_�JE�ZMSSS���U"��3  �D�j6�:88`��A�%��&F����8'Ma���$~�    W�:   �ꅒ�[�I�΂c��aܣ] .��}U�U�j5�J%���)�J�� �X�@�z]�jU�癎yɩ)Yɤ��Y�k:�H���F���Y���$���   ����   \�/J�eI�a:��E���MG0ʉx ��0�h4�h4T(4??�L&c:  #��	b��#��R33�~/@�}rD��c�cga�F�+��L�    &w   ��|L�7Ib?pA��a�\N�bQ�V�t#���|�V<�7;�v[�v[�BA333���  I�뺪V�j4
��t�����
���t"�^��F�#�%}�t   `Qp   �OU�'$�c�AM�ϖ^Z���xooO��7[GE�t:����J%Y�e:  7ζmU�Uʅc �h�^�t\7���c�s��xǾ`غ�O�   L*V�   ���O$}�tDE��E}�Y/� ��z=moo��7����<�3	 �k����VVV����{�1��;��&���c:�Q��y�8��!�a�_��1   �TLp   ��wKzYR�tD�|gKG����w�U�}_�jU�ZM�bQ333�f�� �-�    IDAT�,�~_�ZM�ZM��K�"��$t]�p�~�vԏe��c_0���;�C    ���;   p�ޔ�S�~�tD�|gK-.��`Tԧ��%C5�M5�Me2��̨T*)��� �sG�jU�fSa���'�x��	����3��tďe���D`HC��   L:
�   �����o���� ��Ζ��Գ����T*J/..KK��Y���x�DpG�������fff455�x<n:  ��Z��j��:���8��d�t�b�e:.!�<9;;������UowW�Ύ����������p�)I�M�    &w   �fx��Wҿ���*n�|gK/.J���	�~���믫���=�,�.�^(���y�vww����b��r��|>o:  g���j4��j�x=Q�5�(+�6=O��=�vv�;,���J�Zd߯?J�O�?�`�%���   @Pp   n��$���΁�`��lV&��Ԕ�z�t�������u����z,��+�������J-,({�2�<�x6k -0>�0T��T��T:�V�\V�\��4Q ��m[�z]�VK!�҉8��F%J%�")�}y��Ⱦ�'woO�֖��-�*)LG+��Ʊ/�0O��H�   p(�   7�I���9�A0�<ϓ�J�R�������K�۶���ꜱ-|�T:������2��J--Q~�������J��b������*
 �aG�����܈O����OpONO��0��nW��}����"{��{p@���X���sJ<�����/�   Dw   �fU%�-I?o:���m
�g�,-����cL�ٔ�l���=�(�e���A�}~~8	>Y.K���Āy��^��^�+��hzzZ�R��� �k�8�j���ͦ����o4LG0*}��cͫՆ؏�ݽ=9{{�7���EBja���g�P�n�tDǺ�5   �
�   �����o�����`��mM3��!��E�"��l��lJ_��C�Y���33J���������J��LZDd8����m���\.�\.sr ����?�����Lǁ��=���=���#-�}y��p��Ⱦ�����|�11�2KK�#�$۶9Y7%�`g֎�    @�Pp   ��.�3͘���n�MGI)�GB��K�W^y��D.�ԉ�{rnN��E%�畞�S,�4��>�����@��r*��*�Lu \Z��t:���j�Z
��t$���(Op�,e�y�t
�����JePZ��=���S�Z�(	����#�c^�A�R��   Dw   ���%���>e:&�}gc��x�w:꯯�����������`���|j~~0~fF1�p��t:�t:�,K�BA�rY�|�t, ���<O�fS�ZM�癎����H>�!��$+�6�������^�ȫT�;*���˫T��>�R�Bw&۶MG@4�%���   @Qp   ��1I�"�ݦ�`ru:�{���b���)u�+��j�j5�7z8�+5;;(�/.*Y.+Q.+����Rssx�� �l6�l6�N�U,U.��d �� �n�U��)��!�3^+GI��MG���ɫׇ;`�G���rww���D�ܺe:�H�wn�J�1   �"
�   �9}IU����&Lp?[,�TrzZ����(�&����W^y��x&sj�{jaA�9�������H<Z��S��S�RQ>���Ԕ�Ţ,�2 `��8��jj�Z�}�t���W�b:�Q��^2�B|ۖ{p0(�N^w+��e_~�k:"J/,��0�8��9I��p    �(�    f}Aҧ%}�� �LLp?_zi��{�����Ɔ�g>��畜�Ujn��r�qrvVɩ�N�f۶l�V<��ԔJ���٬�X �k�y�����\�5�.�~�u�)���{�ՒW��*��'J�L`�y�dr��w\3[�w�   Dw   ���I�O$�`:&ӬΗ^\<s�7 I}�V߶�-�[ɤR���%��Y���'��Kp����}U�UU�U%�I�J%��e�R)��  W��}��m5�|���ښ�j�tc��R70�:�v�V���ZM^�2���pB
�Pj~^��L�I��5���5�!   �(c�   0ϑ��$��$V�p�X�;_fi�t����������9��e)Y.'���ӳ�J��)53�x>é1�<������N�U,U.��L&MG \R�J�a���1T���MG0*��sO�5B��֫U��U�*y���JE�Z���Vi�]����p�� ��   Dw   `4���~C҇M�da��|)�q�� �[�>rbf<�VrvVə�gf�����%5;++���Ԙ$�^O�^O�JE�\N�bQSSS��㦣 ���:����Z��� 0	�,)�?�����Zm8e�;|��V*���f�f��H/.��0��k�J�I�]   F�   �/�/J����,���)h0����߿/��}��yN"�S�잚�Urzz8>ux���x�N��N����=��y�J%�EY�e: @��[����|�7���/�W���aTrvV���a���$�����H�Ǳ��1���'%��!    Pp   FIM�G%��� �,��/=?/Y�D�#�����ȹw���$�E%�����L���L���U�\���0�n��n���U(T,���)��
�P�nW�VK�fS�~�t$L���|�t�6�LG ����1/\��%��!    Pp   F˯J�/$}�� �Lp?_,�PjvV����(�S�Z�Z�nl��+�TrzZ�rY�rY�%���}��i���X���$���h4�h4dY�r����Qj�Mj����o�a:�+�a���8�+�K�.I��     (�   ��$���Y�A0�Ǒ�yJ2��L��%
�����Soo�������4��������̌�l���&A0��~Tv/�*�������
�P�NG�v[�FC��(Cm��n:�+`%�J�̘�1�Z����,?-�ߛ   �w   `��H���~�tL�v����i�1FRjiI��M� FB����uy��#���畘�VzffP����ߧ��(��MM)��t�쾳��l6�b��R��D�C� �8A����l��nSjǍ;��?Pgu�t W ����l���$2���H��!    �ƪ   0�~IҷJ�K��`�Qp?[}�׷m�m[ν{�|^"�ޓ����RGS���?ڎJ#�NG{{{��r*
*
J�R�����}xrP��V�#!��z]���M� pE8fq>~��
���]gL    #��;   0����W$�L�Sa���X\�a~k��᧦���^'J%%gf���R�\�oX��m[�mkwwW�TjXv��rL�9�^O�v[�m���(Cӑua��_�E�m�t W$��h:��j�ۦ#`r���?0   ��(�   �k[�'$��� o,��/�b1`�E��V*����SS�&�'��rY�bQ�RI�x���G�뺪V��V��,K�\N�bQ�BA��L� ��v�n��j��y��H�){��_��/���
�8)�\��Y��q�!    ���&   `�}ZҷH�z�A0���~�����DBA�o:
��\W�����&
�A�XT�\L�/����RrjJ�bq0)~jJ�T��O� �n��n��ŔN�U(T,��dL��'�����7۶����H��0�Z�7��M����jU{����x �X����8օ+H�I�A    ���;   0��[�˒�L�xb��|1�Rjq񱓣��~���'�Yɤ������J�ˊ�r�ۉ|^��'�e�b�kN?��0��8rG�JE�TJ�|~x�,�tD 8�єv۶e۶�1	z����NG^��~���m˫���j���ZM�fSa����dn�6adq�W�$�k�!    ���;   0�6$����1�m�-s�6w ��SP�˫��\+�<5�=Q*��OM)Q((^,*q�b1�\���u]�j��t���{.�� ƹ��N�3,�3�O-�Z�[����z]���뇷�VKn�.�ٔ��N`%r9%��uq�u�)�I���    ��;   0����Lҟ7�c�E�G�ܺe:�1x��jU^�z���� _,*^(���;yl�'����~pp�x<�\.7,��R)�D@����m�V��7	#�h��QI��j&��w��fS^�%1e�SJs�⑘���h�c�m:   �G��   ���Z�˒߄Ka������u9Y��^�s�dR�|^��i%�e�s9������\���|^�\N�ryl�����V�5�=�L&�e�|>�x<n8!�I��	�=�eG�o���u����m+8���uy���Ng���s�q���8օ������    ��;   0>6$}\�ϛ����Gc��(	<OA�~�2��L��'
���BA�|~X������'���t��T��U?��S�����p�{2�4��8�@�nW�m�����*Cӱp�~PBo����v[^�9��~j�z�%�{�S� �,&�?Ǻ��V$}�t    C�   /����J��A0>�j�h�[��XL��`���V�W�]�s�������D>\�?|<Y.�ͼ���u]5�A�DbXv�f�J��7��h�}_�nw8��qӑpI���n���~4U��t��>5Y���5<��E���(��	���C�m:   ����   ������fM�x���hV&�����j�t �Q�Ò�X�p
�� _(
�'�]��Aq>����>]�~_�fS�fS�q��h�{&�y��`<��}u:�a��B�hgX>?����O�ԏ������N�tt I�6�h���)I��t    G�   ?;����_3��qy��d2i:���ܹC� ."�o6�?,�_J,�D.'�����﹜'�;�(��\N����*�g���%��Ȳ�������Q�ە�8�t:�<�t��z��ݮ�nWA��~�#����;������`�z�;��h�z��0L� 01b����#�	�$}�t    �C�   O�.�?���M�xh�ۚ��6cd�oݒ��e�1 `���`b�e�Ɵ`%�2�uT�?Q�?*�ݟ)�T��V~vV��i��eşr�<������E��R{@q��ǑT8?����*���Π�~Tj� )��,�'C�O���J���5   �1�;c   `|}��HZ2�������7 ����W��%Y���r��r��ޓ�����lV�lV�Bax;��*^,*����f�����YY�����$�	A �q��;������X�+�r�U��
轞Bו�8��]Wa�7(��z���=x��s�'&�+M�T �+���#ٶ�	p���A�M�    py��    �*�{%��b��`ıu�x �H�I�۪�n�KJiP|?y�+���EY��p�|�PP���BA�\N�a9>Y*�J���dK&���Ǖ(������9Yf?����p��ف��ͻ������t�z
<O�m�.�;��^�tY�u�����Τt �dn�2a��Z-�0>�$��L�    �d(�   ��%��������ߣe��5 `�/�{x9r4�=���y�S�yO<Y�q���V*%+�>��RJ�J���LF�����K�e����s���N+Q*]K~DK��New]W�^O�^奔n�y����*����=oP&?��^����bzx�sN~�ѵ��*d2, ��̝;�#�4�8��I�&i·   &w   `�}����DC�b���Ţ����k*& ��p����,�'58�j�D�ÂŔ(%I�BA��N�����$��%)���JN���5���<*�[�p��L*��n�%&�'������.�;�~o\��u8��v���;8�#�}��=|^��ɒ~��0��:ͦz��^�/Ƕ�t:
�pX|�@���P����NG
�S���W�8�� �f��#q��)I��   ��Qp   �_]ҷK��n�c�1����ܽ+��WM�  ���J��q��d�=�1}Q��)��5��*���aq�AGS���fK�=�X����ʑ8�#p��B�9N������G?�p��e�N�8�:a"�`�wx韸/�U  �E1���8ƅ�I?i:   ��C�   ��F�?����`41���2w�E� pI������cY|Q��E\:]^?Yh  7#9==��g���ǨK��Ĺ�   �أ�   L��J�s���t��/{��� �	�?�<8���q���?q�NG%��$���  0+s���#�!x��!i�t    O�5   `rx�>"��҆�`�Pp�w �$����U~?�X�b7��+������\4  pi
��1.<�oJ�g�C    ��  ���'��;I?a:Fӭ/s���I!; �xT�]:.��u<�=��ǘl��׏.G���S�y% ��b���q��ؒ���C    �:�y    ���I�zI�t��/��*5=-�Z5 �3�����w�k���_�?���m��� �l�;wLGyLp�I�)�n:   ��C�   �<���HzYҔ�,,�]L��]
� ���x���U~?Y���ٻ���������Ԫ�[j��v����$�sI�s2	K��b���f��X*�!Da�:��0a��@0vLX0v �f�m����j9���T�%��ڪ�[���zի��VOKXu���ƛ[��ք��o�sk,�7�ڙ�  $&�oC��wH��u    �E�   �M�K�F�_ZAgXZZR�\V4ʟ��2p��Z���  �\�h]��>�)��W��=�M�o|4,k���:�^gJ�jx�U��^�݋�:  ع��b{�U�
�X�{�n�   ��h6    ����.��t� ��lV����1:� `c�&ϭ���^	�\��p����  @'�3��y�)��QA�s$-[   �|�  ��v��GJ�Y�� �L���&�]d ��A�  ��ąZG�x�|^a��Wѧ�X�w�C    h�N�,   ��[��<I%� �Ǆ��\t��2     h/&�o.��XG@����Y�    Z���   @�����X��=
�s������1     @�I<h��QpǊ㒞-.   �4
�   @x��Sm��8	�5ɋ.��      ��7��H
%�T�Q�     Z��;   ����J:iv8	�5�    @;�����[��xo��[%}�:   �֣�   �%�\\��oqpk(�    �vJ\x��u�������]I��!    �w   ���.�6��A�}k(�    �6J:d�+Pp�kK��-i�:   ����   ��k$�c��I��I\x��h�:     �Ƀ�#t�7��)I�Z�    �>�  ��S��,I9� h/Nn��D?�|�     �O0�}k�з>%��    ڋ�;   П�Yթ7�#�ܺ��/��      �ܷ��}鈤�Y�    �~�  ��u���Y�@�Pp�:&�    �vpA�ā�1���S��I���    h��u     �^(�;�~�8� �ϫ\.+�O�͜�ԧj�c�#Zz��Q��U8rDa�h     t�H2����8tHɃ5p�%r��u�������FIwZ�    `�V   ��U����I�LZ��rڻw�u���S���ОG<bպ��\���������W�P0J     :MtpP��ϯ��/�H�C�4p�E���/�u��㽧��_�4m   �
�    �"�M�^k���d(��RllL��1�<�a��S|    ��D��?p�"{|�~�"{���y�ah�qJա,�:    ;�   H�i8�%�q�1�jL�j����œ'����Zz�������C*�rFI    �v���S��A:�ġC�B��C�[G��L�:�#�t���Z   `��;    �:繒�#i�q�'�/�����k��_���˩x��
G�h��-�<.<���D2     ڮ6�=>>���.R����m    IDAT!%�Ǖ��Bɤu���І���>a   �=
�    j��rI�gA�p2�sD��4p���R�5,�岖��Nz?zTţGU8vL�G����`�    �n�@��1%�?�~�8��(y�r��uDl��}��n�   �3Pp   ��vI�I��:Z�����E�J:��Cڻf�/�T���N{�|P�ǎ�xℊ'O�3�    ��\$��y�)>>^-���WK���J<� ����`hC�[��lIe�     :w    k]'�1�~�:�������b���+>>���=lպ��{� ��w    @�	�Q���;�Ğ<tH�/��8a��3���%�L���    ��   ��,�i��� �.���u��{����ܺ���'%��    ��bgJ�T����b���9gmD����*���!    t
�    ��CI/��!I���!����F�9�}��	���ѣ*;��[��)��    ����٣���W���_��Ptd�::�i���%�z�    :w    ������k���y�v��\,����J<x�:_��t�t}�{y~^���j���	-?n�    �-�XL��1��ǫ����j�}|\�.P00`]�ϴz�iI�K*Z   �y(�   8�WIz��߰��`���E"N~����K���|�v№|P��e��    �v�)~�@��~�@���r���/9g=�ϴzN(�Œ~b   @g��   �\BIWJ����Y�L�B3�Xl�����{��qO�<3���	���%�m�    �,�w��㊍�W'��LaO��+z�yrA`}��{ϙ��q�    :w    �yPҳ%}ZR�8viiiI�JE�H�:
z�s���)66&��/��ڗ�*��Uo�����'N�)��<)��Ap    �/k'��FGSb|\�/T�LZG(����Iz�u    ���;   ���Sқ$��:v�{�\.�={�XGA�s�h}��z|�������Z>q�|��Iy
�    �����J�=>:����
	��9�>�BO8&����A    t��$/�Y`�9�3  ��0-��I�]�إL&C��E"�	��^z�z
�    P�^��6�=1>.�[Gv�vEBt����Kz�:  �l�9�=u6�����D�I ����y  �^ҳ%}K��mSt.�^�i>U��S��)O�T��)�N��>?uJ�S�Tf�   �V|�>���W���طO���S���߿_��1�1���ϲz��%}�:  �|�{���uΕ��1�$ L��  ��1/�Y������'�\(v�y��w��~���ƗJ*��k��q��檏W�����U:uJ�B���   � �~qwtT��������⣣�_p�"�1s9���>#�u�!  @נ������  �  �v����$��:v&��ZG :���W|||�m*���Ǐ�8?�����Ǐ��R�/�8��'�0lcj    �":4T/���Ɣ_�<���ׁM-,,XG������z�P  ������ �{   l߻$=Aҕ�A�}��.24��K/�F3}���ܜ��N�tꔊ�N�x��J�OW��̗ͩJ   ��ۻW��1���Sl�߷O�����\$b�	\���-Iz����A  @W���9�})*i�: sE�   �+]%�%���A�=����b�8���n�K%��Y���|�D}|�$��ɓ�L�   ̹HDё�������QEW����W�HXG���ڤ�oY�   ]�N+��sŨ$ƈ��  v"/�
I_�4b�۰��h�+.��c��4p�nW��T<~\��y���U^�_>v�Z�?uJ�B���  �����|tT���jY}lL��e�����s�Q4`XC�z��[�C  ��D�@&*��;}�{��  �Sߓ�2I����.A��L��!\z�α�/������U^� �T������   :A��_��k(��
�ׁ��gY]�I��  �k�e�@���s�   ��W�/�j� �N
���b���+>>��6�X��S�)�O�������*/.��r_:}�i�   �
��aE��O^��<n\߷O.��
�E���uNI�\Ҳu  е�}�9G��$~  �ݻF�#%=�:6G��m.W������sn�K%��Y���U����W�'�ðM�  �/�CC����QE��_)�Gk����S�LZG`la�S�]�"���~b  t/�����[@_��/D%�[`�	�  �	J��.�ے�g�&�٬���!���X�:�rlL��Η�*g2�"|�˩4?��J	�V�/�<I   g�����퓋D���Lp�*���)�  ��A0ｷ���B�{�R���Z   =�I/��7���Ypa*��jdd�:
�.�ѭ��P充3S�W
��充�D�LFa�Զ�   ؽH"Q���g�b{�*:6��޽��ۧ�=g���8���(�w�;$��:  �~��c� �;��!������  ���)I��������)�h*[*�K�/�T�fם
_Yy\���>^X���
  ���}FG:�xp���A� ���ҒJ|I��'�ْ�  ���!�6}�h��� �oι�3  ���&I���	t���E:t�:�>�je�m��+�|u�ܜʵ��\}yinN��E�0l�{   �Dѡ!EGG����QE���<�����\|@�[XX����-J�\�� @S�e �A&����	�  ��^$�$=�86���t��2|r_̩M���r�"|y~^�l���\N�S�T)��   v.���NR_)�G��_��)>:Z/���V z�au�P�K$��u  �;�0|(� y��Rl�D�Zg   =�(�钾!�|�,Xӯ ��Zl+*��J*/.��ɨ�ɨ�r_�d�������E
�  `עCC����o������E��>_YU�LZG S����pno���  �������u ��sG��\r���QR�:��s�寻��zի��  ���SUK�wJJg��l�: ��*28(]x��Y;!>l�_��S%�����r*-,H\= ���8]=:4T��VdpPѡ�U֣{��E"ֱ��Pp�h��4m  ��뮻����lN�֦� �5�l6{$z�WV�������u" ����s�3�  �U�*�zIa�1� vf;�%ɗJ�I���p�_��S%�[��<7�r>��w   ֳ��RllL���Ue�h�r�Y�����d�#`}�I�B� @�9�|:����_���ĿNOO������s��;Ї�s?��   zޭ�-�*� 8��� �.����ƶ�O���J6����٬ʙ̙����a>_-�g�
�y�\� �u�������aE������ޏ�PV����� �rI|�  Z�����HRT��s?���J��� �v�Zҿ��k�AP��A �\A"� �P���F���+S����Y�++��Tjѻ `g6-����^[��/� :�au�Pҋ%��u  ���}��io��n��	��  ڤ$�i��t�8��A �E;�_C9 �
�� ��gX���>j  �X `�6��Vp�w�?�a�]�  �oU�ҵ_�4`���qr Ш���|�z_(����J>��PPX(���T]�˩R((\Z�$ (:8�``@���"��)20�������Y���\,f�  = ��XG��K��  ���� �����Rp�t�a v|,��:  �+ߐt���I�[��r��*��"��u @��M9��W*��{>_-��J����*���2|��r>��Ғ�ʶ�|^�� ���j�|`@.�P$����P�L�.���Ճd��6+� �	�#�껒�o  �H$rO�R��2�w���=R�:�>&�Y" m眻rr�g�s  ���vI�X��w7�|����k ��
��d�����Ҽ_^�����׶����+����"ey ������x�\$�
�zY=H&I$��j)=����I&:�>�~G  4��^/zы��u�~wRң$��:  �/�t�~I[� �>��SSS�3�%�^I�m	��=Wo   V^%�%=�:H?[\\�� �9A2� �lʱ|���X�����j9�P�J�z��R,V'�
���R��_�X]���P��T��@�H�^(b�j�<���bՂy2)�U�I+� ���W{��W9�� ��r��v{EI��v  `�Qp��s�;�Ǎ�{D��+ι{�3  ��Jz��oJ�y�,}kqq�:  ��b��b������%)U�����j1�\VX,*\^�.[ZR�
W�=��Ru��6a�$_((�T��?�o�,��,I*�r-y����䜂DB.��F$�s��E"�y4Z/��h��.��}�x����F��@��� @��+s^իp~�:  �Oι{���Y� �V�Nk�����s�& a~�:  �k�&�+�F���%N `�V�mU�~=�����\�/��Pa>/I���aX�4�+U
��~��佼���l/��~e�f�0�>,���3�K%I���W
�>���b1�$�)�K�Ҹ�j9���ʿ�ιU�>G�����A��A+�DV&���\<.9��ʱ�����Ū�^  �>�2w���b  �/��7�3 h�z��^p�F�_�pY\���a��  @߻W�%}DR`���p� ��S+G�sl��T�����p�eE���:ˤ�R����S*�R,n{�F.Qd�%�`�~��DB���.�P��^�֋��}k�r  ���d�#���$]o  ��H$�5:�@����x���t:���ڞ����R���  ��M�n��o���+���      ���������Y��G?��(I���   �����{�u mq<�J�_{�jB�s�i�@���u   ���t�u�~�,      t*>�21/�2Qn  �{O��_m|����8�@o���  �I��+%}�:H?Y\\��       ���{ە$=O�?[  ���
��U�ֵ�/�7 +��/Zg   X#/�ɒ��/(�     �S-,,XG�'^�u�*�  ��A@��ι/6>_Up��rߐD��}����=�!   ��SIOW����     �N�gWmuXҭ�!   ��d2ߑt�:����ݸ`U�}zz�,鮶F`������:  ��.�E����2�      �T|v�6wH��  ������s h�/^}�ե���-��_h_ �s�� �N�aIo������J���      m����[�3%y�    �@��}g���Up�D"�2 z\�R��:  ����X��u�l�:      ���^�\�:F�{@ғ%��   �K�tZ��Y�ֳ
��J��v`�7�p���C   lы%}�:D/[XX��       ���d��u�^� �2IY  ��J��>� Z�9w���_�Ok��Up_qG�� 0���u  �m(Jz���X�U�L�:      ����u�^V��<I�X  ؆OX �2��knTp�У�s�| �ns\�S$qV�8Y     �N�gV-�%�J�'��   lGtހU�T���^����f�N�G�^t:��~�:  ��#�
U'���8Y     �N�gV-�vI�X�   خ�.���%������d�K�X��>==]����F`����u  ����?Pu��daa�:      �
���[I�[�   ؉+���"�S�9 4ݧ������V�[p�$��_�. ι�a�  `��-�u�^B�      ��Ϭ��^I�I  ]�{O��=vZ7,�g2�;$�W#�;Ng2��[�   h�)Im�W0      ���{S������A   vcϞ=��t�:��Y�`�+3lXp���.x�?ޚL ��{�����u  �&�#�k�Az����u      `
�M���TIZ  ح����$���������VnXp��H$���`��g  �c��.�t�u�n��B      t�:�eU��m  �Y��t���qΟ�s�?/�XS� ������/[�   h�9IO��ەL&#�u      ���6�J��   ͔����S� v�X6��¹68g�}zz�,�}M�����uzz:��  �ߗt��/[�s�P�L�:      P��U�v���u  �f[����:��q��������Yp_9�{$1��^�s��S  ���%�L_�ۡ���      �$)�˩T*Y��fwH��:  @�8��-�b���y���f�lZp����Oҗ���ϥR��X�   h�H��ѭ(�     �S,..ZG�f�(�b  �a���?u�}�:����)�J��f�mZp��S�t!~~ @9,�ϬCt#
�      �|V�c�I�}I�    ��!�8�Km�ӺՂ��%��U" �d2�  �F���:D��!      :�U��IO�t�:  @;�r��Iz�:�m;�G���
�K�޹�H ��9w���t�:  @��D�g�CtN     �S,..ZG�6�Nn��u  �vY����u �㽿u����-�%)���$��@�X��6�   ʒ�!�[�A��ѣG577�r�l      }*C�������M
�~z�u   ��,��P�D"����n;G���y�s�y���ݜs�MNN��:  ���%}U��Y�&�x\������p���e���S$��     �W*�4??���y���i~~^�\�e
��:n7)Kz���X  ��N�o��R� ����T�[�8��#G"���aH��|�9��   ƎIz��%���t�b���Ǐ����n�Q~hhHCCC���ݻW�m�;�      �@�RI�\nUI=��Ջ��|^�lV���:u�*��u�^�%M�r;  �sA�=×h�Þ�_o������N�ӟS�$�s}"�J=�:  @��UIwJ�c���b1kppP���;�_+ɏ��)����     ���zc9}mq=��)��knn�:.�7H�c�   � �NBғ�s 8�ϥR��������aRp:�s���   :�ݒ�%�c���Y�V�T��ܜ���t�ȑM�_;~m1���      �MYo����y����0�����KQn  ����aRp:���Î ���wy�s'�h-��g'''�:  @z���K
����b��FFF422��{�jxxX������p}Y���Ȉ"��ul     �-	�P�lV�L�~[���l~~^�LF�R�:6Z�IO��7   ����J��9 �뫩T�7��ӎ�����O�d_ ����	  ��}P�!Io���*�J:}��N�>��}�񸆆�488X�_�_�5N�߳g����F     ���h�z�V[����癰����LQn  8KoÐ�;Ё�0�ӝ��k����J�����%�.�J=�:  @��Y�X�@����ke�Z9��߸|�޽rn�v    �.P+��������/..�R�X�F��O�c$��  Щ�����o��*_K�R��Ɏ;��.Ia��];�@�y���:  @�F�IWXAw)�*����ӏ��-�S+�ixx���񃃃��S�    ��ڲz6�������z��9�J%���}G$=Q��  6s��W��d�!�s;���9�N������1 4�GS��3�C   t����Jz�u�Q<��𰆇��g����hdd����|dd�>9>�LZ�    ��,//+��)��*��iqqQ�LF�LF�l�~[XX�/+�ֱ���U���    �`vv�����Y�  y��vjj겝��	���a���`7��kIl  ��%=Iҗ%���Y��b��ӧO������/�kttT����&�7ޘ    �F�MU����eLVG+Hz�(�  lY�\��H$�d�`�� ^����L������s���q �s�=���/��  Ѕ.��}G�1  �IDAT5I?k�0A1    �.Ձm)Kz���X  �6�����޿�:�ϼ��}jj���9Ʈ����F"��I�� �H&��  ��QI���$���Y��+�:~���?��}�Ѩ���544�꾱�QQ>����     Z�\.�K�k��ճ�l���:�e^�u��  �#�H����3%����%�ܮ��KM��.I�t�5�^ߌcضT*���  ��%���C�������V��Q�   �&��4�����yy����O%M[�   �f���)���u�9�^399���g��%)����H��f��}?��l  �|S���4h��Y�bQ�bQsss��w+��������    ��YA�\e�b�h���$��   �6<<��L&�I��u���(��4e`sS&�KR:��\���:�-��T*�)�   =�ɪ^��6,�c6+��b�U�4�Q$�~    z�z�R��j�FS�k��9�Iz�u  �^133�D���s ��{����Ǜq���%)�NR�e�<&��y��zjj��9   z�s%�OmV uk�XL�D⬩���c���\S?�   `h�	�[�XT�\^UP_XXP��o@g�KI/�  �kfff>�{�u�OܑJ��Ԭ�E�u I*�˯�F��$i���p��H$r�u  ��I{%ݬ&)@�*�*��������hT�������@��xK&�J&�g=P2�l�   �O�P�ߖ���������jϗ���%��햖�����n�t�u  �^��s�	�Ƭ� =.罿��lzYcff�Z��ۚ}\ gx�_>55u�u  ��jIo� �'���q�b����׶i�&�F��GFF�p�
   t����R��b�x���b�x�T������|>�L&�r�l�V ��g%=Iߜ  h�t:�rI����kS��;�y��ܧ������������c���_J�R�w�y�,   }�m��� �V+����z9�V����������
�   ��4�΋Ţ���b��rz���Xd_XXP��o ��+��(�`  ��y������$��u�G��%�\�W^ye��mz�]�>��0h��~��Kz����}�Y   �Ȼ%��: t�x<�d2�d2���!%���Z)>�Lj``@�dR�DB�DBCCC���J$�u�d��<  ��R����e---iiiI���*���rZ^^���
�B}������
���Ţ�����.--�X,Z�% �Tߖ�XI�    �`vv�%}�{?h��1�A�����w�}���%ivvv�{?۪���9�����[�s   ��@�G$=�: �x<^�_�$�ŔH$���k��'��b1+���  �Wզ�7N;/���k�����޸_�9 ���Q��>o  �����WH��:�c&R�ԟ���-+�OOO��ß��V��O�s�����]眷�  Ї��>&�2�  ��i,��&ȯ7E~``@�H�>y>�ippP�hT�DB�dR�ht�z  ��h,���e
-//�\.+����/--�\.o8=�X,�P(�*� ��}�~K�1�    ��{�fgg?!��M��r&�y���tؒ��5�>��=����u�>p2�<����:  @�K����[ t�Zѽv�v�|�4�Ƣ��}�N���bP�o ��q�I�R�����q*�z�k�d2��e� ��K�͕{   ���9���W��,@�[(���馛Z��MK�433���Z�:@�{F*���u   (!鳪NY ���ɤ"�ȪR�����Ѩ��䪩���d�^�w�ippPAԏU+�מ'�I�	 ��
��*��
���0���Ҫ��|^�{---�T*�P(������B}2zc1�v,  �ਪ�)~�:  @�K��O����9�n�����[�-/�KR:��M�K��Z@zG*���:   �%�)���A  h����7>n�H��6����ݯV� t����k�����Y���N9�h������=^ZZR����  ��iIO���    ����}�����9�n䜻mrr��~�h�_@����5��ÿ*��x=��|#�OY�   �*YI�#�K�~�8  MQ+�r����f��J��488(�ܪ)���%ihhH��D�H$$�>�c �D�·$��yI�O$����eU*I�����ƥ3�Ͻ����Z2_{  v,#�2Qn  �(����L�W%��u��ܛ�d^Վj�wI:|��	��nI{���@����?rjj���A   ���$}Yҿ�  v�6U�9�n~``�R}�|߸>HZ]�_��_�p/UK�ιUy� �?����N��]S�T�pI�ޯ*�׶]�,�X&�M��kiiIҙ/�ݿq}c��{�J�R/� ��������  �����o�$�~K�� 6����T*�/�x���%iff�J���h��]�{�655�q�    8������:  �/�E���������U%�D"�H$R�v�}$���kje�����x�F�S�%����Z����&�o$�������^�X�>�B��0Ϲ�\.o����V��]�����Xk��a֋ݍ�X��1����k���s�(j�r  �6[��4I��  �����<�9w������gMMM��v�`�(����$������snzrr�O�s   `K~N�)L���   �}�2Um�   }�(�Y�n�  �����L;���:�ɜso���|u;_3�|���f�$��~]�[8�n���x�u   lُ$�����   �}�Ţr��9o��  �NI�D�  �k�R�?��W�9�N����_���~ݶܧ���J��\I������w�0|�s�o�)   :ȏ$=N��     �~U��BQ�  �*�9�U��oZg:пT*�g]y啕v��k�ּ��o�� �.i�U������R��X  �����/I:d      @�����  ��I��?#�$�o��'�0��n��/��	�5+o��%�2 ��9�w�]N�  ���P�c%�      �-(�  ���e���Y���{�U�]2,�KR*���s�Y�ʖ9 c%��3&''�n   M�CI�%w      ��Qn  �!�T�n��S%�� �*��799�U��wI��������9 #�{���ħ��   ��~�j��A�       Z�$�E��  �S�����bI�:`�{��T*�Q��wI�����{�z����LMM��:   Z��+J�      @����?h�   -�J�> �5�9�v�޿~jj�f���4J��o�t�u�������&�s   ��~A�%4�      `�(�  �t:�FI������R�ԫ�C�tT��{�fggo��
�,@+9��>99y�u   ���$�)�u       ;V�t��X  @{0���9������9�u���:@#真��|�s�6�,@�׉�����   �⻒� �u       ;R�v  ��399y���V�@�/�ɼ����R�ܥj���/��$��:���f��-   �M��~�:      �m)Kz�(�  ����r���N�,@���K.y���thd-g`#�{7;;�g����4�-����Pn  �{�"��ƭ�       ��v   �{���t�97a�h���r��+:��.up�]���g$MZgv�9����ɛ�s   �cPr      :�v   �233s�s���9�]���́u�sq��T*���:�,�y���)�  `�{%=Q�	�        �U�t�(�  �����[����Ա�``�K�R���r������ξ�{�.IQ�,�U$�"�J��    �XWu��~�        �j���n   �ivv���wK�Yg��✻frr�V� [�5wI���}��y��� ��y�������A   ��(�      �#�t��w[  @g���y�s�%��l� ���T�#�A���
�t���W�T>���l�����SSS_�  ���I�%w      �RIҋ��v   l��Ç��'%�o���iIOM�Rod;� �511���_��]�,�:���?�r;   ��ے#��       @�*Jz�(�  `&&&�Y�T%�n�,�:�T*��r�ԅ�kn��ᥥ��K��:���x���^{�u   t����I?c      �#Iϒ�q�    �N333C���{�u`ŧ���o��� ;ѵwI�޻t:�'ιת����wν5�ɼzzz:�  ��w��%�_�      􁼤+%�a   �m��z�s�?K
��9�ޞ�d���NkO��ggg��޿[��,�;�J�R�  ���_Ւ�í�       =,#驒��:   zG:��\�{%�ZgA�Ytνtrr���Av�'
��ַ��� �����:��s�[�J��n���Y   Г�I���GZ      zТ�'K��:   zϛ���K���_I�5�,�ߓtE*���u�f�K �p���f���{�u��;��=�v   ��iI����       @�9%�E�   -r�M7���G�m��l6��^)�K=4������s�s���;��N;���^�|   �FR��H��A      �pR���m�    ����Wx�ߩ�U��f����������4[O�%ivv�b���$=�:z��+��U7�x��A   �w�n��{�A      �.���'J����   ���������r�=�.�΂���H$��믿�G�AZ�g��w���/s����~�:�V�{?���f���C�0   �[QI�t�u      ��H�$��:   �S��*鰤!�<�Z���?��NkO�k>��0o����Y�]�s_.��/����?   :���IWY      ��wU��~�:   𖷼嗢��m��ߴ΂�� ^611�]� ��wi�7_ҒF�w{�#WY�a�y�lw4ݖh��J
H �!�"	�E�`P	��L��"d0 m�j�����e�ƽHJA�!����B�@����s^?̖�B-��3;�/��O�yv3�d��yO�ս7��v�����I�$5� �\�:D�$I�$Ij k�3�7R�H�$I��Coo��1�>��{T�Bo�y��3ft���WS������t���
��OC_Mݢ�B�]�R��9u�$I��7 פ��$I�$I���j�`g�I�$�}���N�1�c�z�է���j��ŋoJ�2��n�[WW��B����-�υ���啩C$I���t=p-M��N�$I�$I� ����C$I��������cS��n�B�~�\�e�
�RY�j�?�̙sKkk����@1u���c��X,����X�:F�$I�VS;}��K�$I�$I��� J"I�$�U�Vm8���>88�:07�M+��V��;w�hɒ%Oݓ�������M�7�,u��M��Z�^�hѢ�S�H�$I�ap3M�%fI�$I�$i�/�� 1q�$I��O�-[��B�p#p1������BW���SǤ���]����*���S4�	!,,��Ϥ�$I�F�%�π���$I�$IR
X,N"I�$�����c������N��wb{$�pU�\~:uH���>z{{O��|)0+u�Fݟ�<_|�UW=�:D�$Igw�S�H�$I�$I�(ݩC$I��Ѷ|��,[
���E���,��J��R���{���}
��OO���Bx<��e���H�"I�$�����O��$I�$I��� ppG�I�$i,�lZ�n��ٽi]�p�!����9p��)4��7��:;;M�"I�$�������C$I�$I��1�� x8u�$I�4^zzz����v�ow��Ú��/������<� ��{�v��ʲ��\.?�:F�$IJ�j��;&u�$I�$I�4^�6��[�I�$)������y� �pPLݣ4�̲��T*=�:�Q8p����ӆ��.!\��G��B�}xx�'�-z)u�$I�T�����$I�$I�F�������C$I��Ժ���B����G��B��.��/��i4��Coo�G�<� ��"�=S�����b�����J$I�$ՙ"p�Ӭ$I�$I��F�8x%u�$I�TOV�XQܵk��!�K��pӚB�ܚe�ݥR���A���(Y�|�Q�B�1�K�i�{���!�;B��J��R�H�$Iu���8u�$I�$I���B� ���$I��YOOϡy��Ͳ�{1��R�4�7��Y���T*�K38pe�M�6ͦ6�05q�D��}�q�ԩS�7o�P� I�$��� \�:B�$I�$I��.S�H�$I��R�dmmmsB���n�(Bo��1��u�9pC�J�#S�L9;�x�`J��&� ������ϟ�+u�$I�����B�I�$I�$i/�\
�C$I��F�bŊ����Y�o>p�ہCwm߾��J����A��qR�TZ���f�.���{�x(�xo�X|�Q�$I�4�����!�$I�$I�D�F���!�$I�D200Pشi���91�s��S7ձ��6�+ݴ��tuu�B8�p*�}��6�1���;;;��:H�$Ijg@[�I�$I�$�}T��"u�$I�4�uuu}�6�$NJi;�ݴ�MԌ�ׁJ��2y�䓀�B��Y�A���ҫ!���y��zƌO���WSGI�$IM����L���$I�$Ij<o��N"I�$5�����ƍON˲lv���'Sw�����1�'��;w�\S�T�SG5;�u���o����,�N�1|80u�>�
��1�!<U(����x!u�$I��w<��C�$I�$I����M"I�$������j�:;�xb��� �׀gB��<_����dGGǆ�Q�_�H__��CCC�gYvpp��u0)a��B�q}�e��y�>��lKK��lI�%I�$i�<�:D�$I�$IM�e�,`m�I�$I{���?mxx���qY�����!�#���zӺX<�����I�&����x%a�>�@�Riikk�B����4`za�[B |l���:��`ʻ~�v`�mvQ�f��#�7�m1�W��!��b�[����3gnnoo���)I�$ilM� �N"I�$I�����<�:D�$IҾ(lذaz�P�B�c<8(�p0�ݴN�G���M� �-���#�Wc�[��Y�m�1nޱc��J�2�� uG��\�    IEND�B`�PK
     ���Z���  �  /   images/a5640015-ff5c-4848-bb8b-6d4b42e5489b.png�PNG

   IHDR   d   ,   ��U   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  eIDATx�՜{��U�����nw�����n[����Db(����!J�Mj�$`$��	j�/�HH��"�JA+[JHw�ew�m�5�;3~?w~w��tvf��-z���������y�o��з�?��m���G�� 7Z0���,�HX2�������0s�k`�����gL��b1�f����㑑����6444�f�qM&��cL�7��Dr��vy�ZKK����Y}}��������'��sm����� �(q�	�@�N�b��z q>PH#�T�����q__������?�u��	��O��&��-�¿袋�q�TKK�1	fX�Rz`�Fzz,%��RB\+�Vs���ga�#i�C�ʈ��}P�C7�ߊ��=��`	>œ&M�z�~��u��z��s�9b�<�=z���L������Dr�x��R+M@ )	s������^�A����n#���֪�I�R}0�c�l�P��r��S����J�0�N��@��9Ӫg̰�E��a�76� b���p�4���O���������_�y�B\'��MҤ��->y�%Ĭ�Vw�V?�;&��9��2��i� �H��wX�=">t��4�'-Huu9�<�S�[�}�;���c�ſ�'�ZXQ�7�+�0��!i���n3W����N���&����jC�����[l�YgYV��0+��  �=�����G�3�/�o}b����s�lD L�D�|�����\&4�<@��Y.:��EHQ�P|S�A�8ٙ�c���o��2��>�Z���A��Д)6 �����>���H��ng�`K�);?"��-h>��
��O}�x���$-h��얦�459-�;�d�|�IϮ��a����Q�+*�E�-���Y}8rV$&#!�'$��r�PeK�Xϛoھ��[--�K��Z�T�='�O��0m���6�	�n�<;�3�i�
�1]2Yh^\��u�0@�͞]HC P�U�E����C�+
��dav�@���6[~�A����6._n��l�SW�����Fנ
 v�{�HpI	�J�̀��(�i��i�P��ò�������NZ��� Ǥ��ɣ� "�el� ].���e������4��T���g͝kS��q�B�u��G��S�G�Q�'?i�n�����oC��oq>C+��3���f������a]��u<��(-҄�{�؈�cQ0"=�Ƣ�Ծ"��"�� i_:�I7Y	���Y2U���r���@�*;팸V�k8o) � 14�A�(��ߨ�5��A��t qy ��,]Ӧ��BCF�8>���9>`�� �����|"�G �`B�	>DH|c��Z���1��@V�X�����6,�&���p�*g�d֪,L���߽��B�O=ՙ(2����Y�;DB��X�@�"�� �;Iya�e�D�:=Q�V��p�d��ciiW����O?�&�U��d�;}_���f�\�L >�4M�%= �)h(c,Ah�� '����Z�ż�je�Ah��� �B
�Ci�7�~��,sW�� ��*�Qڂ��g�~����8�|�����SOS���.���[�mVA��3����Ѐu)EM�.��������޴�!�iO�򓆏ܚ���<�'���=0�Lr+��g���6N=�D�7��_Jj}�U�*W]~�'l���g��Qѝ�h�RI%:r�t���$p�������euO���]�I��Y�0xH�*����KQji�����x�&]3Yf�Gt 5�i�\E�J�mmc��ʕ+[�j�U���$>W��1����K/ھ}��:�O�3=_��de����R7�U*�]I����-3C����P~��m�Bט�V|���u�F��b�sk)6R-�)��B����1Ν��޽{��r�9s�g/�䒃ZhI{o�:�ϋ�9�%u����t{�0LҚ5k�D��/��PEݣ�QNw!i���  ��LBP��@RҞ��Id�Z�Iq"(s�DP�|�r��瞳9k׎�'�@l�Q��o�V4֯�1��ء����~��2�oY���������2���+1(6|�+����}�'�
�g�����Kve<�Ջ��w�H���,%���.S��1�FM���_�+�H;b�2/cb<z~��EΌƂ�� 1��˗��/���XF P�P08�$�k �yk��U42R�J��g�e�m[N�EV�c����D��G>��d_.g��-�K/v�Tň�1��^{�R0�xo�] Yl" �bb
�Q�!�wA����Bo�A�s�Ǜ��@l89ߔgr�#��^V�/sc�̵��{����TN ��wK����S%4�
6�<az��\�U_�u	$f�>P�U4��b�	Y=Ŵd�sD3ʸ�V�@�ԡ7�d�?��")@I46�ayb�i���DdUDK�[�'�HT6����|��n׮]�lٲ�N��e��%i��֦o����U��͒3��o�!q9�r�(��b;vX���j
 0G�Z������R�(*1W=�����7���q*���EN�LJhU��e�y�66��{�Զ?��+� ({ �I��ͽ�Z��<"SdQ���/�}()A'�*�2ǃ��H� ���M�M��%�r yD|��h��I�s�9�7�|�o�k6m�d\pA��p�:_�c�z��R�B�4]�S�|�8܅�ҹe��\~yY������h��ڂl��~��kL-B3H�������>�쫷n�ZN��fϯ-�f�K� �
�*u+��+�D����k��?�p��ɵ�]g�Ѵk���e01��2x�%�F�DZ�(���=�i���g�7n̕��!%Bj�sؕ�b��������y���u_:��Γ@yiݺu��\s��I%��@F��o�����B�'���l/�7EV�|rɞO����$h��K����Ü�~�V����My8t˅����wu]��v��YR.�za��(�j�?,�Q�a��ʝ�ehE�D6Y�A/����-�A��4r6���ݮ۵t9�U+���c����z�Jd龺�-@��B�\�@J�5�_�
S�t��*��x VnB��z%�&�0�����&sqP~ �nݚ;nc��;gv\7#�p����T���Bh�pM�g�� �*2+D�l��j�p����a�#��+��;��i�v>��l���4c��EPhBF;�ۦ�D^5���ٮ�|��E#,r�-��r����m��	M�d�E@Q򨘢R��*"-V2N��cr�����ޯ�P�7s�jg��?|���`r�#�	�K,`�*��lL�������=�a����i0�����������$b�|>1�l��7bss�[��Z���7��d�Ιc�
�iX`˷���`��Q {-��^�����BX��}o�aIi���뭍����(�8�'�����/���g9γ2�l��Y"D�S��̟o�
����5b{�g��Wd���C_sN^��5��hM����|W!�n	SV����:��6�����G��H��l�+^��ɲ*!ПECB�݌!%_-�ۙ��cG^y����uM�԰X�'�\��#��a�V|�|KMk��+D}g�v�l�fS����~�1p�؊h�,��E(����Y�%hL/��#�z��L{٘���e�}J��D5�]k�2M��6[����C���fk^��E:߭듛7k�l����9GF!3c`,ɠ_��@n$��mQ
,j@v[�}�;��zI �n���Ӝ�p@��A	�[��0�ޜ�f�r�k���HؽA���@ �o�n2>�W��xj��/ �d�@��"��x?�4���s�&K]�� h��x�YǾI�s���3v�h��ӵt�Pv���]f)�c'I�\I�p�_槏r(��O�$�ڰKI�7y��aB�]�?, ��[�T �w�{�%�M�e�L�daR��"�=$a�g�#�� �3�\c�@��X!�ہ�Ycc@�+m�sh�hX��<ely>�l�ާ,J�@���E�)YX,�x��������l^����%ָt�h�@�:׃(	A��nE��������$AnłHilp�����'De����x�>c��O���q�z^^��+�~a)Y�I��\�g���ſDCz�!׽A%տME�W��;��"$ڄX�$w���R՚��1���;��(<�G#�9���1�Կj�{�/r�Q ��x�xi�~*�b�#���klx��Ɯ@�������?����z���|9�8����0ή�R��9��V��� d��-�h�'D��x�����{9t��r�1���x�Ȓ'����Ev���,'_@�g���1�����b>8 ��D    IEND�B`�PK
     ���Z	��} } /   images/bbfae99c-8036-4c5e-89fd-a87441410720.png�PNG

   IHDR  �  �   ��ߊ   gAMA  ���a    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD      �C�   	pHYs     ��   tIME�#Պ�  � IDATx���{�m[���Ƙs����8��GսU���袍�i�4��A�("�q�6'9�Dq��E�HEVd��HX�d���&�Н��g=��n�}����ךs��?Ɯs����{����f�J������k�5�x��p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8��}�𵂪 ʳwQʄRZ����k��{�Lǁ�%O�h	*T�J�`011@��#�QD
*B)�@ FI�"4"L�Db4��L[�>T	
4AU0����11��*��J���N�L� ��m��l@�(`\m.@aW��7W�G�|������%���<�Ç?���p8��h��@K�J���s�H��K���EFi��_j��R�kh�,A	P@	`   �jQb���!f(PA�U{�B8��W? � �FE}E��z�T�0b��P�t�>��1�yPr�P)[��7���I�����>P�+��T�hT ��ۻL���J��ui� ��5%Nd?#��z�vH
U�w�[��}��rV)R�""�%' ��f�v�U!�bs�!lJ���x�/.��Σ�~�S�����G����7 xD������%b~�]  A�=��~l�,!	"bz���
�*�E �
$S�
t�Nb�Z�L�WaEM����DՀ�Ĭ
�h�AU���!7�(���?��˯���1(��a��%�۽�����]���$���}i8���U�5�ժ��T�[T�GE�C-�J��eC�����	d�VE�RM��F���dQ�liO~M�?'0�w^d^�b�Op�x<��L�$����3x� T"��q���/@%B���w���w��ڄ����k��3o������k�q����:Eӯӳ� e�n|�Z��	U�M"�7h�Yr��((W���� D��@U�����y��䟽��� �6� ���X��D%"H�T�(�R��0+���	|KLO�x��8L����m.��>��m.@aa�]�%����P��/  �Sm/�J��eM�7h.�SD��J�$_+t�RM��
 ن^X�f��@�aJ��QS�t��k��纽o>c8y�l�BqĻx<������{MH��sF����J�v�������U�v�+��K�������]^\��^��������ԟ��|�^�/�-�p����; t�0�>]=����_.���FD�[%���P�)	R
b�K)PUÀq� ̦���2���_�+t�;������2{��W�~N�D�DF���k��q( �fB8�g���90��2�d�����q��o}a�X	�@�>�G�ᗍ�VU����n�./��'�����/%�n���Z�K*%��Pɦ�T d�ά��H��Du�Z�9��yeӕ�����}N�]�v�W-�~��;?��c|���	s)(���QJA�fB�C`036�`6q��F��,��j�@�.�q�}�_o��v�y�~���g��W~Ƌ��Ǉ��q�`ڿ�_�o~��-������<�Β�o�o��V�|����D2��\!���!F\]_#�(Q�W�Y7ƽ˧3]oqǕ�\`S���"ZM"�� J�jTM1+���y����M`��P���ϙ�gƟ��~�Ke�q�1^\!��1��,���;�������/b�]�����U��HI�Z2 ��"	���`^yۨ�j���l&��mH:��@��l�
^P]���u�{	@��9��s��{<��s�7��.���L@��i��%c��؍6���1b�<b�#��E�0�+l����U�_�������b|�_n���7^^���, "���~����g~�G_�2��W����O�����%�v��7�i��|8n��[���R@*��PJC��`�!9���E��^z�U쮯�(��RU����� p� )�z�5���5ki_2����&�5���5�Ye.1WEO�����9
�'����e~������3������1ݾ��}�������o����!����?��9�.��T��9���I�"')�
�慢�B{�g�Z{�^IU��mt�Y�8��ieٮ����$��qԮ�0Q���.~a�9|*���ÌL���9�((#cF�P��BDĆFly����.�<`Ѐ�p��Kx��|}��[����/�~���T�O@)������W�������~�ǿ��y��/a�yʘ��b�]���o�Ͼ��2r�~��p��3,����4�P) ./v�$ bLsƓ�^z��x�ʫ��
� "���ӅA<�t����<���])U��kH��Wy��P��]��� �r��G��C�U�/J?�!�(��#���,o�M���#���#��p}�����u�П���|�G�|���������e��_�|+��*�Z��BHU��(t�ͧg}	yK���*3
�U](y%@hM߯��@���a�y��`��s����N_�8�@IAA���`F �!�b�
��1�6<"P t�J@���p�勏��W�`xTv���8?I<��ƿ�H���4��.��C   �7��+��4�i�p�x�xx<D
�:�ߖ�߭i��A��8o���� � �3��Md�H���#��9g�./����g�N	�^~��������Č@=Q�z�I��;:_���LV6�^�l��H���_׾6	�<vQ q�P��@���Y���q�� �o�D7x�c����@�P���/�*��A_�����폐����_�^�����Ayz�� � �J�h�V���c��S�w�Vν~I5!�)t�j�/%]š� 뤸��P���x=@B"��%Ct��@Q2��j�H1�Z��JI#2fd8!% `@�� 	!d��������F��:��?����R/�t�{C�o���6=~��v��o�~�qw����AU�RP��Bd�p�:s)�ó�?V4��9�ߍi���p��·m)�I��{H:@JB �%�'H�(iF>�Q�H4(�>�@cA�	�M7�i��;()D �%oz����q�9t�:W�dg�o�;��#����u��I�%�X�a���|����(�߮y�#!���@o}���8~vs���[_�N
��~$�}�y��޲,� �Q*��9�%��kXӀ2A҄��4�z�P���oYY����aJ�E�*��j_�*�cYXk�PN��l-(/4;��.�S*7����S�����	��IZ
� H�H�.� K-��"
5�d0�6؅+\�x�W.���xix	�0"`Ѡa��4���g���e��2���x��p����-!����n��K�u����9��3 �����͗���o�*2��O�\~_��o���O�i��N��y"�3Ho�Z 2!�#JN`"��9!��r�0�nn )!��8D��r��E@q���5~�۰���FFV3#R0Yc���Q�.DW��ޛĉ�~��P3	j��6��*s{ͪ���O�u�y�T�����UM�0(�X
�'a:��C�i�ݏ�{|����Ȓp������/	_W��/}�!l>���(�Z��-��D'@Dg�(D$��I�\��%�-h�Ӿ_|�U�v7Zy��1o��B������״}��;��"�ܴMȋ�iT�b B$�j�,�JBT�[J�A�X���B� �غ �H ��`@)B�6(��3o��4��4 �	�kL�c�O��g���8�0��s�Ͱ�~i������w1lw��t-����@��m�$�9���M<|囯5��۫W?6�~�j���K���U��n�O!�-�dYfhI�r��-E��	I,^.9!oq�y
��0n�u����3�4�c��ͣ�-bܘ�#��a�K�J��J�S���$�U�ng9��޳�R_T�9�h�EƂ�@�����OՒ�J�I9D����)㯕0��D�ߺ�<�����~������������O|�ʬ����O�ւ�Z��!�㿡e�(�)G�r�j2[���T�<s��qن�R�T;�Ψ*t���F��9��z�Z&'銢jT�4*���-���9��ւ�Y�]D@PD
�H%�&����Q�VC��H*�b�#Ka�]"�Lϰ��pF��~ʀ(
�y�&��M��7s���Y���t��1�� ~!����g_�t�3�C ¸�Ї��43�3���/�ٳ=��
WWeh���u0����#��̀�rP@b-}�j%A���BH�L@mX����D���Iָ���Z�X�K���jZ����1�}��p�b��`@IJ�A��AT0� Ί�2f�vD���q����Q��0E�t�c���
����v���}����;�y�%��j`���A����o��I_�"��>z=ݾ��*�E�'E��Z�5D8���h�C��	�@��|DIGS� H.ȹ@0�	ДQ�#�t � C���05���uw��"_? �&[T$K||�7�ӄ@������u�{��KoΏ9\����%/D��=����f_tN��;EJ�֛R7J_#�@uF)�e��{�O�����~����~�w~�w�����V���u��o��|���W�|��K�H���"G�L�2�lJ�%ͫn��1F��Ϊ
��w�yL��M����E)��z�ž6^O�:��׾�aU �Z"@�lB��;��,O�@����z!�$(J��ށ ���l���p0R�Ť���3bQ\L��-�����A� ��RB�v������5���������3S��8��"z�oso!�o�?�O?���q(1��%��f�tv"�w��T�Բk�a � J�s�a�q���	L#�iF�G�M3�:Z2r���<�������}��ʟ���G�q���D��2LE��FG�b�c`��B���L��	, )�M��`bb��Y��I ��H�tr��7�>½�
�����_R�U�Fji����P��
U"����V!�K��R]
E� n�b#��:�Ah�t�����p!P �����^������ 8>y��h
n�S� xh+�Q
�60C�~a�.�J�s�JB��g�o��}�f�g��]4b��� )�����/�9^
�Hy@�!��H�q���7��oW�߂r|]U^*%_�f�P�W�Vb�%��@�y�e>"�(ǣy���-e���'@b��%c:� D�4�e����!�@nn��gL9B9X)Z) ��oN��%�T��G�ÛR&��!��Xe�$��nғ�A+��.R�m�e���Ξ-�K��%�i3 c)lT�D@��H��)�''�o.����nz���O��#���a_+|���f-�a�0o����5_)�R�Ũ'�H-+SA˃T]�oQ�a���g�8M�X�jU�X�6ֹ-���s��2�kѩ
Z)�wR��G�؅["D�Ь(�0A� 6A�(g(B��g��#B�dU*`Q����)^C�
�hA��43��A�!��A�^�^"���{�BxF����D�%����ox� �q����ՌF��� r�0��N����N3�W��z���y `_��"����.
D>����d�"ø9��IidC�qP�AJ� �1�C��n�	1��R؍X�S�4A ��(TsE��*7�\5s���C��L꒮oZP�7�7T�/IAbJ]�i*UΩ�Y�(DETUE��Q��q��THJ	�E��,Y@9�EU���PJ�&*��"���T�\��-�˂�-Ƃq,�~�_�9�B�R����٫Z��*���l��r�^�3=��C�<�������`�hH�޽P�E�#��HyՇy��\i�;���9�ΐ־Y�'ת
J� �(%[-�<��#��M	�fS�R ()4%d�ӌ4O��0#猔R�P#�b�R��0����f�� sg8툩9�M�5[���Kύ& ���K�{}��$ԭ����ԍ�ƪ��ηváv�_=]��p�b� �d�I�oU%��w�VDE�n��2��ܼ�i\����zV��*�ӻ�'{�q�M���/i�sH�G(gh��V�V2���>���@��L�QSƴl�N�t^~��۷}JQ{]/1��Q�&�v���^N� ���M^[�f��FR�`l8��#v�E�2CHl�Q��I�d���I�zp�`��DDe	 &&��Tn��u�b@s���\KE2�L��  03�Ja$#��� V�P�C��8&���(4�(QS&��L���U���(I��+���� ����k����v
�<;��T�i�����a���2���(��r�BsR��H�L��HDL̡*_��i`Bd!��͆i�/]1^}i
�U�K��q�u�V�����û��|Խ�6L+MD$���Ｔ}L_՚����R/n�7o+%Y6qVe) e0���([�DDC9BDTPP�([P�P	[`���P���VG��"�%�HI��R��Ǵ���V�!T�T�c֜7�������Z�̌�{5Z�v<UHUI�����V��b��*K� RX�0����b^}�P�*��g��S�Ħ�i�q	e>�oQ��d�Ϥ-�Rl��������
���cJ8���%��ْ�b b4�:M{H� �S�-iM�@cS���YS���3=]<4e�L��&��7��D]Q�2<f-��w�n.�~��G5�,"�mb%S� ����Cx5���k���n��4r�x��O��Z����~��C\~��雟�m�������'PI֛Xg@��=��F"�j��V��w~" O��~M��S4����z�}�,���歯�f͆��ڇ�d��fc5/{TƆ��BϬPeX�2��Q�D��p���� +#h@�!����!?E. �ƂѕD���huRTC��� �"�z��`G�� ��o�����Z�&�Qz�w��y��CUf�<eL���O�xrTd,�X2B����$b�:
�xf�<�3{�D*}K1�ĀAB���0!h��̀a�������D!�����жt����M޻��o�[}����F�,��'����ͻć��ď*A���Rt�-^V��$��%b�p��[HA<a�`� ���tܢ�K��щ�P��-!l*1AF��lbM����l�=Y���
{?�x�=Y��k�
h1o��Ĭυ4�C(�"E���T{OT�ԩf])tj��u{#I���|����) �֬�~��j��|D"R��<�8���8D���M�l"B$��ʼ� ��7S�(�i>�϶լ^�n�ﲹ�l]���{��*���F��* �:�et�볰<+2O�b芚���ĕ(�Q	Py���P��}������ȳ�O��)<x�[�aǇV��~����@���4���n��*�
��5Ͻy�B���4��*���{����z73׍ghq������K������������E1[���
2�P��  ���
��b,�F:� E�Rz�A+0p(��\`��y
(]Yk5����C#��jV��!�׃V�q���#�g*w�ξ(�/pW�j���1�$I @�3n�7�`�@����D�;WDP�@T0�	%[�b)&l+8�b76RT�	��U�h�\�	~'��}����N�25�6��~��	Z�"�	"]��l�
�{��)T��!@��t��i��#Xf��`�
@cy��4@C��-hs�v�n�p�{_�U=4�¼(��8�2�M�[S�XN?�m�(s�5	x.�5>�3��j�I�z�K���O�,=f�{���'��=@5�\�]q�P�#����JNV]R�0��V�V�3BP�t�����^_B&3��R�t ������ߢ��h��t%��2�O����T��^/�k �Tma��0�����?{�J�KM�CϷ��r�若�E�� ������������'���{�	�|�Sx��oy�g���R��޾�gሇ�UM���K:��G�̖"�f�Ve^�~	��!7�l�n[��%�ӂ�-J����ן�)z�+��O7�J�wLZ{Rj���5�X���ʜ �2�H
��N
S�\@�M�Aњ�7Ȥ"(�}ge5�t�@��r�1�A��`�8T��湒V:��}�*�%j�ΐ�E���m�"H���:��`�ύjڽ���D[̀�� �#O�,RD�l1gV�@��5r.�sF))���!R�e�0�-."a`���UjhדX�3���=(*x>V���-LY��u�� ��=�u4� pT&�NвM7
SX��0���vL3(O�<�'j���J�TD  <��:o �%�`�ov ���^rZ�U��Ր�5-mMZ�ЪL�p��Mq��g�n��[Bz��֥��m�h͏��_H}F�Xy�-��׽�O�}��)��a��$	��L77fP��
�����mă�s��2w�v�n��Q&���	6�U�!��o�N�Jj�u5��]�r���5[��ht�ʘj\���AlD���^�Q�2�~�*��~`�L3�j�Q���`���69W`{��$
�����O�G�+����`��e|X�S�
���ޔ|�'$�T�<hIF�kF��PG��r�V�V�̓v.+ֶ�Im���'V���wS�k�ܳ[�u�z�<��/[�]ey�)��ԪI�l���w&�v�@m��d0g(�*��%����6�%P�Q����4`�r�$3����л���ٵ��^&*�W�*ШUi��P�,lM�����Oj��w��(W�kJc�͆ ���Cf�"(U�81B��� �\��{�V0P�Zl��-×a��|Ļ���u��
H��O��T�C��]�rQ�͋�=����v��(��b�.�`���.��9�ƺrD��L��Ϫ	(
� �	�� %�����T "0,��T�2�)��!� V�._�� ���M�	b��GX6�+��:ٻ��5m�*��Z7�6���S�|��β(������h�Z={ċqQ=z�RKK�2��,Dl}�I��,N���9�!0(0r��b��#f�-V"I���`I��7�f���ۍ�<�?`:$�3dN����z��
�:٫��{�����5��x�M�wơ1w"+�[��`�G�����\�3���}4̌��OU�#֌�z�a	J�������9=���G���'�����q��gq�!m@�S�7��T���%����%�XӒ�e��l-=�]����+���f�����j��$��Ic�٬R:�컀&+D�F�¼��,����*�C5Fd@i�DA����2�b�'�f5+�Փ-( R$�FիoP��(2�5��Q��/#c/��2n�G�A���vo����Rf�;2\@� ���l�r�@�Ӣś����O�\ʲ2wj���k=1�B�l@R0b�u��	9<�f(P�le�2Z�p$F(&���d����Lur�Ֆ�R��
�12�����x0(X'�&�-���.���[����J	P�o�Jm�tU�띪�ꋵQz��-g�R�N_Dd���	:�V#���Wg��
��`L�,IrU�TD���*
���n!�-�b��PF 5�����B���O#�-�e	^�@lFT���<'�6N�5׵Z�ֈ��贌����3�L�Z�ZmHͣ�&�+����o�
o��vT((�e!OG�)a�8B�`�7�W�����O�<��֔��|�s�LG��"6q�V�K����YyY�nJ����^��:��*p���T���85�~�4�3�<�ET_������J *5�*˥�v3���k�$9�/!��O����ç�K/�>T
}z�H��'�|�Ki>|���:!�)	��lJڒF�4�Tzh���Bk1�"[�R��tE�uO��V+�����oS�M6,}�[}d}��x��
��!PH=�k%�����(��`�)�X��>6�	!��MHP��D	3� �z�,G� ݮ����,c�f-�|q�5�u*���m�cB��5���+/H� �������Ѽ��x-$R�9�T���9�Br�� 8��ԗ	`A���
)3�
���2z��@�R���RlT-�R0� S��`?r��y�]>�k���ݵߴ=q�e6�Z���<�~��{j��mˡV���Ȧ�+���6*����D���̥� %�L�3�c�j�V��?GS�f`�	 {!*��C@k¤�A��^I2&��0)jߘ�%le�w2�K�C<�<볳ؿ���[;�K<[����V���.��*!��m+��Y0�*aD
D[WHE)���h��!"�3?~�9M�\I�a`!������./���/DH�1����iF�%3�焠-n^�U(��Da��O7_Ջ���׶6'������ڴ��pL��idJ��.o��oK�]�����M��`�Ř��>��9zB� ��o�7_��v����[��/�>����Q誊��/!�Ã��͟+����<�J2�\l�o+�`�D¢Z�E� 5~��$�d�F�-�k�}+v]�D7VX2�W^�J�T����i{�	�槣�!U2�bk��Z'��`�[v��kw�~�%2� n�>�{�8ҌIf$(PM�#�f0pD�4� &�����܎$t��Q^)iՓ�5������Z�t�i�a=�R�P.��	�2$)����<!���JѶ��1FcD@�hID)�T��"P��{�Rޥ*-�K�=�z������(�^�VN��BJ�F�<�u��'5�AD�O���[�q[y{FEP������PB������ws�fԁ��B$���0K56YH� P��8��1�8�ᵕAB�~i��s^���^'���w��DO�ZU��_�.��B^����!��?tf�����0*~=DJ%�>���Ŝ��[�yBN	77Oq�&�֫���k��/�q��BDPR��`���'����'8�(s��4M� ��j�����@M�yW������BS��o���3�(���Bn����\������nșaѪs �_Z��%�ތ\�1�������O��;�����]|v�o5�&|(����������9������<�ђ[R�1b��%�Y\1KY-~�g�7ũ?���@��y��Q�%�ף�(zvh���3!��n�;�@�����7b�線�F���J�Lv�"@z�0{�v@Ĕe��$�P�g5�V"w(3&9b�	%�`W�}��j�����#@JFN�QJ�`��P��r �լ����h�"�(�F�׷�>k��F��Z%�2 �)f��~5\��@�i&���y�R�#�1 F�u����"�!�keA�sQ�T�Ů?FFL� �ϧ�q'˵�H盡��]��8`�ce���4�e��1&K�9��
϶΀e��ʘ��a�:im�|ʼP�T��R7��{U�x ��h� T�ʆ�5T�/D@f�<IP	�o�������c)��%~�i�n�/K��C��nG�V`(j������k�gM�=�S���I�Z:o�v�TK�<"BQ��������equ��d�>}�y*H�#R�8�v�ǓgO��l0������)%��<�\
�	����Gf��%l���7u�,,�%�ô$�َ'9K�@�r����:�җ�3Q��6�h5Z�:;-����)z�LY�u�2]�r=� ��2�������Q��|y���ǃ�+>,����"����]|�o��S����<}ea6��՚��I
�-~���Xr1�doz~d�z���������j-a�3�W��X��L�L��1*#��e���5_]p��aM�5�A{G&�L`����Q2a�#2f�Z
 B�� ;$��5�02�x��F��x����0F�U����W��r�%	���,KZ�v���߮�sk�c	�F�.��j��S�-	�Z7S��pn}�T�JAI�s.AB�H� �(IPf+�4`�ڎA�%F����m��J�5o�HWR��{�'�����e�`�t��S^�g���JʟP��fL'��d��`��ք�Z��e��["�P5LXZ�F��s�X�n{E������9ke+��u�v�1��Q^+�sZ:A��.9�gJ�mW��E�����]��wj���/	5����p���J�Q����R�tx�iNl//��G^�~������ FJO�1��r��a�ʌ�xDJ	Zex�)�sO}���a]���㥯�k�;"��Ȩ��\^c��V��$����z�S�W����I�z�^#3$��6B���?���/������}��O��cߌ>p��������7�v�돤��?U���J:�%�D!ɐ�{2��R��s��r�~��K&o#�j�2 �z-6Ӕ���9x�ڼ�x�h���z�,����|�r-be(b����q,��2n�P��0}��S��j�6���%aFƬ3�L�2c���l�!�pG�C�ц�l ��xF�R���,�z!��OX])t�$����x�,�{_�V��1w�J�
��� �1a@ҌP
B�Z��X )c.Y3rJ��>�gD�F���E)+R*`hQ�ڞ�4�*������S_���5��[h�y��������0+����e"��Q�EiA��iz�7&2Mlg�$��0��T#+t���Ĭ-�ь 5�Ό.!K�5�l�n.�����ڪ�_)�x�ٛAsj ��v��
���F��I�7���W�S_��("]�o���9\Փ�����QE�d�C q@*�<g�R.8'l6#�FpQ�qy}��|�u���x�����}�� �i�8L38D[����	i^�,����3��s���Qp�F��$c���oxnI���J�\�{j5�:+��8n=1L�����\�e ��L	N��
I>�����0=}��}o���x�o��T���%���ax���(��G�|T&�Z��6�	4Z��K?�Lړ��k��S�Qd�� K���Xka���Xv�2?��Kq��/8��V�t��=ʿ%C�6��"F���������ѫޓ�:oAT�X�M��Fւ$3�L]�[�j��z�bε�e�vW���8>@���:C9#�Yp�����S6���εRWt��}�L��n��lb1�w `�)،f�
��֖��c{(KY�KR��X�%�eA��`�C�hQxUkKlԟ�n�?m��
��;Վr���G-�g�hԽ�h�*���! %,^��>FcQ�GҌ[��5-�7�޲��%���q�8�&�ڡ�@�Pڹm
�Ң���[(Gc+Dj��T���E�:/����K�����װ��Y{R�H���3��(��#pzx{�W���2o�C7ԛ���3*�[�@ss@�qq�4g\]]���#���8N3�d#T_{�%�~�d)x��cd���T0�qs{���{�a
��rFN�ĠYd��lRks��t���8Y�;����K���:�������H#���ۺ�I�Z���~���B[�f	�"��A(vn�:m?rI b��t�^��/��>���;�>��ۿ|`
]U������_���{~����h>��2A$�g#����	�j<]!@� �Z��&&�-�D;�5i:��d�V�D�P������e��k���y�H�b:������;�[Љ
;�Ӈ:�KA1��0b[�Q��)����ژT�@�2*�n�aP����lY�(�R$HP䈩�"˄P�B	�C�Ad��$A�%=����!�xe�j�!<d�Bt���&a�1)���u��{+���E��qq���ŦTJ�BEj��"�pE�����焒	4bX:X��Ա�@$BΊTj�
� I	b`��`?�΄cV0�d=�j��P�h�0�e:��I��v% +ͣ�̖��R
��.���?ۗllPh	�U�	`LK)(Z :!ȡ6	1!�4����$"����JMk_]�F&k-j]�
��l����������4�����	����E�֑ �)YIT��ֹ'���ւ����v�m[v�,�Ѣc"]�-L�:�gevF~�>5�n�Y��+;��i�����w�l/����ݣ+l6�4�����f��^������	�b��<���,'�x8����r�m�{5M���#'
�}y���vΔ�q����L���g'���t9 �o�u]����C뫯'��Z~�U�؜�j�$��I~�������������߂����|�o�-�������=���I���t� 5���,Ѥ��-q2B�Y�u�A��ن�W]j��.�`��O(������W5��w�Z���|�$윾�Y��\� ���7}A���[�U-.W։)�M�b���,����f9X'�b���-CY��?:���@��:C���L��E��������� $�Z�o����,ٺ
�nNUa��ߝ%�����D�c�E���m$"d�q��fQ2�T�p HY�&�D"D��`���5z*�\�X7-����o=S<>�K대dzZ�*ζ:XNH�ԖF��=��c��Z9���a��\�Jw�)Ag��^"E! J1_�,fK����rWB����Lw��(�Evk76Hm?��[	(��a����e�`�|v�������a�Ӄ�&�E�5�Q��f��J. �}�j� h�H�S�f8�Q��q����z�-sga�Z�jkKZR��i\ (6�t6`ETPJF�'����#����a�-B���RJ��v��	2�9c�#a�ݠd`;��n�SB��)8��)M�P%�J�!�,,sKe��{�x>I�<Y�;G�����z���c��3���Fw�c/_���>
����:�	l���a.�24-�D"�%A�d��_���y�}+�>�<.}>0�>=~��똏��W��GJ:��Ɇ���#���T�]J��Z��5�^��K�.ٱ���ߟv�[���`
y�1�f�)�=v}rg_��(],����p
�u� m�.�bD`
��jrגd�(�H�ſ�P���EfZj�U�u���Z�EY��U�	a�#�	*���H�,�ea������DKM�Z���0Е!Ж��0�H(�\=j�GV@R��j�s�&��J�zܘ�$"g˼�LP@����Aр���@V�����L���18��ߺ�qCN�����CS>��;���@Kz����q��ǵ�U ���mF�V�3C�2їw_�Gv^�a}�hM;��Ty���"���d"Y�Bɦ���-=y���=�P��� ��"+O�5�i}�W�\=c�)�O�w�V���*I֝�t�m?\��f1�g��i��[_��&@5A���^�j� ˄i>b�#�`�MeZ.���߁����A�f3"��'X�RPJ�dWǨRs�Ob�f��f��}u�V�ק�)�ޟ��q�峽�����Ým��xr�r"_t]]�Ƽ
 *���=.�2�1���O�g���?|�����	�������UzH4g�o�B��$�w�:9M{)Z������dP9��E���U��Xj?������[��7�*rfMU���ݤ����sZ�Z2%���0%�Ɇ���&�B7Nl���i$��5��דs��SR˜O��:#�D��#����<�;ͳ5��d�&�N�������`j�nBAd�z��^/�s�B*�lXw[k�o����[���L�o�m��a� �%�Υ�Bd����T���U��CR׮������x��w��?���Q�]� �����s��vJe�X������֙��������J�+b�!��i��[+�:e��#v-���K^Rm���/�ql�^�:U�
ъ�4/{CZ��v����7BNAulks�AK|v	�-�	�>9�X��*��_���-�R\
3n��|#����)��A�@ ������vLs�������^sr��@���%��n�#�<M�ӌ� ��<�w��u��{KM}ϟ�����-���'��:z�*���V�ja=TÔ5�Xȥ�L�Kӌ m��@Hy�.�����|��o���>�m��'�s5�Z��+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs����|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�f:���E�s�.�L����)������@��w��{n�<��D�^K6�md�c�pcs��yN���I]�$�����i�!�����9�x��=���b��ko@�[��E�S��y�a1�F�bf���W|��	�64졻V�#���޵_���d���є\[���0�h��9N�	���N�!�2�}���2c��?�ߝ��
���{��HI��z$��W}����7S��o=�|ֶ�����]b4�3R. f$ʠ̠\@egJ��%�Ȼ=�T�4�h��]�8T7�1�j�{ȷ#�i���f^���=�d�w=ܲ
	�1Hg�|_��O�Zb#��cE-cm����>AXj��T M�Z�iF��3ي{o�GE�z�E�8c�v�7�n�6��e��I-����#qs��F{J��w`f,�y+ �׽S��=Ӵ���Í�����WV��H7h�!�kO��6վT�#��N�l�N�E��O�2��e9~-�����!�xS�U�׾�19��?W��NH�w�ȥ�"��x{a�p����Zĺn���|r�j������!,}��}cu��o�2�T�6�;�n���1tKY�&�!{��1��]�}zߺ�F��t�*���ER;�H�t����ǯ����z��d�a��x��iW��Hcx��-`�*c�&�b�ns�z$�o�g�{/E$\#>����ЅQ��HIM����+$'�4AZ2O~� ��yM]#�ߌxn���%���L�ځ��ہ�̣��c @�b^�l��1.��cch��}=��&4��ƒD+oB�#��G=t�b��O�Jid�m������>uʫ��C��i�&�T+n%+n圁��){4���g�$��J��kB����ͥ��V�ƃ;�:�J]]w��{�X�?�:�&���=��������O�m�j���*V�����*C�=,�!���*č{��UD��������ݣ��q�=M�\���58.ɚw�iY{���tG����U�-��~���7�O�o~�e���� �il0�C��Ъ��m-r�� {�sB*;P�~�S���� ����x��:П}�{���9 ���r~+��H�X��ԭ4���}�o�@j�#]�^�*$ [KR+�#��W���s�Ƭqtݱ��m�|�6�]�ݲ$�|zYh[=�=��{zQ���f`�{CX��]cX=
�եz�e��i* 5�¾Ag"$����LDA}L����vA��!�Vo��t�2vۤ�o����j���ĭ>�s�����Jk��\,fqO:5+�Y@�����`�083L��&1���e0+r��guU(ߚ=�/��N(d1���WG�1!� �wX��̽���z�ͷ�kߓ�XQ�d�:x����I�H#W޽Y#)���:M̢���t�܈+�$K�d�f�]��D&I^�h9��� M٢>�w-���ugQ��������[�˼`�ŵ��ͫ��}{{���F?n����%��m�4����>��	�s귕��WHպt K���S����TPe��Ċ�#�ہ�Z3!g��tlW}k�Մ,�c��xh^Dp��Hy�Ϙ�)\ER-Z'	@�>Q�ڣ5↳�BU��?��7�������a����^{3D��m#�2ڂ\�������$"�w��;��9�8A�
��r��\ (�N`ڻQ[@y��Ȼ?��?�7�����?�7Ձ �����_�9,K��n�JOr��ip��0���P��NԚ�x!ء�:*K{���G�������c����_���pc����YĲ	k�Yi�L��M�0i�>�O7�77������ɼ,�l{H�7�Q�L�F&��5ܷ�R��0�> �c}����5�%��� 6���m8�/�Nv�j�$~	��A]<a�:s#\WEU=������hJ��-R��y�x>�Ɋ���p�4N���*�f�kǆ��q�'�:G˩E⑏��5�QJ��E��k;������0<�/tv�ֲ�"�PuHޓ��i�l�����'���f�71�:�^��)!!�Y�F�i��^��̮�X.���R�.��*VX^�6�Zl�^X��t�Ϭ�$C}r�n�I-��g�����]��^�W����X�����ӫ\k`�f
p̌R\��>�4�h�v�UR��5ۏjkX*0�Z{V6�͕dG� �_�{���P�u9�I��E���5r3��#�Q���-b7�"]���=j�Q�d��^6��SF*djp�<d�X�4y�������t����w�Agq�����~��K���7~���NzE~�HY���h2�7���rZ=��a�]�o�2�����,k���m�cV9�߬�'76Y�hm.pϫ��Pݶ*�o`�y>���r��e%�y�͐t%� �V�:B�6�I|��9#�y���@N	3^T}x��i; ų�ÓD����5�{�!�l��彘,�^$�)2Ī�uV�M�M� r[<�A�J��`��ŕK������J������@�N	�^��
4��Sww��3�^[/���ӄ=�8��I���Z�:�����������>+�X�����:�^�u[���՝t�+�48�b�/��	>�N���SO�)�&9�5�~h+e0'��m��R�C1��ٌͨ0���z��A��g�y��������@"t��q���z�7�\\��Ū��Vḧ́�ך�_l{�=�$�ު���j\�J���r7������f`8@�V�	)OÐ�V��d3�ن�����u]�P<m)^i,zlp]��v��{Iלޮ�n�l��gA�m+���Kߺt��"������ϻ<��2��	x% R�(�<�ly#�I=�)!BJ�א��s����2�^���A��xS� P���o{���?��~�����|K%��M~W�̓���0��F�Эƞ�j��e{�����@�l��l����]e<�}'H.[�19{xh�gW�z_���
�0�y1��؄�Z�W�ZG����f.���X7��X3#b҂ H�$s�x�i&{���3k��!^?K�ٔi��@���u���:�6a��#^6�x[�sU y�V`n ��y�P������h��=�f���\�b���m��	˲@!�rBNdS����̣*��|�K��]$�W�����f׍y�z�c�S&�������خ_���[���ӱ��f=�����}� aW��e1/�<$��{�잒��!�Ecm�׾�\���@+�2��<	��$���,�v_�쨧��K�6�MX�/����ֵ�][�_;����@�/k�}���~��x�ǟ��vcٌ�_����o�=K e��6�~Y��� MpCI��n͢�Sbp���^Y,(@"F���ڈ��LP�H �)��M�3�،G�{(6?\1�q[�G�H��U�p��9ҿ�h�����8�8��=j�w����!�c��E� W��8O�#�8'(gP��T�<�R�0=��~2��+ǫ{�=���Q�y����~��﨟�9�����Ͽ��?�����"G4,X����C���IA ��۵J�ԇ���R�^/���O�6w��鮘�mB�:�D-�	�.�V>�sQ�Jzh+���R�2]�!�ILloߋglZP?_��IU��b��EO*�����t �4r��mU�g�{}�ȉ�h۞���?��26�5f�!Cү
�MR�Q�Rd�3��n��{���K2V�,��V\^6<)�L��Vۨ�ruh�S �U�d�3 ���խg�!e3D̨i,:��յ���޻�cܧ�g���ՙ��z�F�9��SztC��9z����~���M�A ͞̳�1r�������WkU�|4e@���zw�}-[�;�-���}
��]�2�Ț 9����ģX�0���y�\�|���q�����#i��n?-g��=6�k=��n�z��X��kU���4��"�%'L�	9%;�`�L
挤�T9	@�l�Fk�4r��CY��
z���M�B܈�\�H٣~�������zQ�p��������7�����zU�Yn����n���zU���{�*m�ל���@��(Д�����7�\��mJ{ ����ɟh��}���aqޤ�it"�~����Ư��q�����OO	��1�H��֦�^A����e�B�aH����#T�k�]M���C�7��ƚ�G��.[WF�yzŪ=�ݳ{�_�(Z��Z�V��Y�_���'Q�VJ�D��Z����3�0��t�6v�����"����)ﯕ֜��ٕ�n�9n����X�g�W�ۡ�s�.w+�:Q�M��s���e��+\���-S�n�qy!x��@� R=�n��j/SL)#1#�Aa�2RS�g��L4[;���抔3���L�\@<�6����h��q2���zR�b���M�j�7����Gd���{�CZe�EٚK6.b�֘�(2sF��BW[ߍ�
2�L�T��y���!����sF+tqt�.��y��@/�Z��wz�Q<�]O���zM����Y@���U6��d�{�Q�p��l�x3 s:o�!o����{�Z��li��~�4M`2�k��b�dbO�JV1�'�ͧ�l�*���*cؑ�v9EWEi���O���Q5�e��`|@�����ݯ�*�D7��X�vO��,cF�f�z=Ł�ߏܻ/w.�^�z:]�L}w6c���{p��yO{����0s��e������ `�(~���ެ�it CB�s�(�|]./~��<x����0��ݽ�q�k7�M!��湨����z��u������X���æ�lv�&44���%��t�9��#��4<�ѿO�屛��L�������y�Խi �40��v��`$O(��K��;�m�%v��IM>��=3*(�9�++	�������ٟ{� �:Q�W�JU���QEէn	�������Z�
hJ�1-G\��oy�Ɗ��ZQ[C�L���PB.�zf��y����&X��V@����ē`i���PJ��eƝ�~���W��&�9�f�mk�p�)*�zlN{t	MҪ7��w�Ev������aHٌoej���v;�a�r�l:�P�6��&���N;H���A@*;�i�@��'s�tq	=��.�8����Ji�n��a3�'7�ӣo�`$�\9��#���l���#2�kH�+���p�ѝ��Þ+��I�^���}�Wd��[=���m���b��n����N>��B�x��-��V/n�����G�9m���\�\zAl�
jd����å�>i�H�!��G��,����U~�������H�)Rqs�~�	�ŏk�EG�f��;@��kDJ��C��Ɣ����2퐦�T&�r���i�������S�����7���M�M}�w����s�(>����������K*�	Q����˧���9���e�ՕP��=r`�ʔ,TBCAZ�^�Yվ S?�W�����z�h-�R�ԳC
O���Gچ�\�]�F�����Ⱦ �(�a��B��@�)���j���[�	9�0Q�!gܚv��.pQ�8�=&-��9!��vJ�>'�Z��ۃ��d�ѣ��MW�z���am�{# *r�P�̌&�|D�'���l��{��	g���A����V.�Z��ǓU�i��3�
�Q���a���	mO(��e^���b��dnD*NMq���'2���t+cAc=�t1��}3|��^�E���t�Ve�*���E�x��;��}^wJ}F��NH��9���=\��&{b��кN�y<�i�`KM`�ВВ��!*�߃�'!w��g0JbdΞN�ϚR�y�<��7d��(�ի����U�&��[����Nڣ?�Ag uY0��=?SA��K��郡l*[�N�
�� M7��6�<��#�,H�L�`ڡ���&�,�V�'IR�tEj{��p<][$*O�i�z��CS,�tid�r;��?�z�9���"M�������[Ov�)�S�Z��E�v��6y�.��3aҸX#�}��+Fl_�}��
'���#�����-��:X��D�+�?��2A��\,���`���:�>ޖk��G����S�7�o��C�3�0n������^~��9ܯi��+𣤺K������|�%՞�@nM{ۅ􇗺����V����V�@�W��X���K��m����xo9a��Dmآ�E���ƿ�W;���	9��5�o]�@2#%�BJ�����[�`���T�����3i�e������%v(v%SvO P����=����U��>%�BA���H�_o�̬Tv�DBDJ�oӴS����'䴳��4�ݑ[���Z��¢�V�dJzJl=����`�k(�C��&�s<����&03��Ќ�)�J.���-|�Kh�Q���D6��� �	�+�d��'2�'�����б�������Ƴ�j����ѾǤ;����/xލa߽)����?�+T��n#]6�\lP���*H:���(B"�5���R&P�x�M�4�����m*����S�˧�r@&'�V��o&���5ZU��`���Ƭ AM�A�H9�%e&eb]�E[�*M�*n����������N|�����M�D���'�UIDIUHd�Jċܴ��}��.��0�X�R�)_�̱��� ��?y;��3)Ӕ��_@�p�X�()�	cވ�Z_����dެx�@�!���RaKM�}��M$��IU��u5�!d�(�5�;F��(���F��7������7�S'=`�=#��h��SA�%���r�;�:��ns�3���j�������\��|Ͽ�����?1�2: ����_�ٟ��˸������{�=��$���酪���k��+���q�����f�KI���ja\/"���zC8b�=4z��r{@������G����xiKtE'�zPTm85A�#�d�c����>)I�"��gMH�(^�iyfFJJ9`��\pk���t�|�|@!k� '$0)Zv�>�����������S#JU�-��DG"����> ½�t���!�'�{<pՓ�^K[qF������
9��*�*�T�lҞiwU���v��}-�:�'ngpR�Xt�@p�GiIN��2��e�t\x8N[D��v�D�����E#B*��pk���-­���.����yL��X r��k�ivD�2���MWA���vf����^�E���Y�U@�!��. d*����
��Ҿ��4%�\4��!�"������3v���O@�L��K��'�O�佧��̤��&�ĩ1s#BUEm�.�<SJs���r:��� >NJ�>щ���隠G �rﵓ��"h'-j�,`���W��(���p��C�])�n�����>�|	�U=�&��-mr)��փjۋ�I[+R[��L��$���"�T��HZPX�XG�\���).��)��@�KL��Φ�ժh�J��Ac�>TB����H��nl,��&P����=� �
�V�Aɮ��;�ױH����}���I5��u�g���)#�؝��*S�g���X�H��{��}�E)�K��7��v~��,�Q���w�9���G?���
~���=�f��˷ԁ ������+��q���_hy����m���<1��k�/Q�"%ki�&Hb�0i�N�:���*&X�ܛ��x=��hxI8������V7�U�C&`l �U`Q�PSA&��V�'�W ~�0)R�P�ȔL�L2�0�f1QA��r��i�;�ܙ�`���<!���VA[`�ښ��Y����T���<�Ӄ������5f�� }�2^d�<����h͉+���ݾ*s��n���ҔX.�����2��r��Sʍ�y.Rk���&�eB]
8=U�߯����wcW���������T�E�ITx�j���P�'n)�4/x���Ǚ�JΦ���	9eH3)K&����S�>+n���pkG�mFW"D���+����}��6̨��m�.o�J]ꛣ�^�lm�Ex���~��Z�.���. �Z�����	uf�(�H�V��݄S�q:	��)���gԚ���%��ٕJ�n/|�����S��#_3�Cb<,�����_�į xE��,*ߨN/��[.��[ޕ�)7�,�rc��D¹4"m��kd�e�&Mx7)�De�k�,�jEz�Qr��m�@��r}dL�y*iJ�K�Xu�mn	@Zj˵�,�%�9Km���V淋���R���|�H}mym~B��Vkˡ-ׅuIB�mAʌ�����q��i�����B�N��]ɸ�`\��КE2
d)�vB����hb:]��HPP]Еۈ H��u�Ż+]�����dE�"����Q�;��'�#u�BDS�;oM�{爌Z�q&�a>�@0{�>���>xe�R�#O{�2]q�-�������������R�9�-x�v���Ox���_�{��Oѯ�ҿ���A^�E�� -&�)&<Cb櫶il��R����D��dZ��\���lz�{��f����!���&N��@2AQA3�넂v���z�����+de
��M�1MH�=�N9{�3�JW�c���].pw�w����z*C9!��Ҥ�,Dt��&ί���Μ��S�\N�O	��*��9O'N��ʇ%]ޞ?�3?]�|��r��R3���֟Ih�J���n(������-���Vlr�js�L��'���������9\\�5��Y�q}��YQ�KD�[k���i>��c��[A*Y/��P8=��J��e��yλ]�23@���5��ä�ĉh_wD�/3������?����²]KοNە�9���D�`P���F�1Е�[�pV(�GE�B��:V��� �MՆt:i�_B�	����Δ���K�Zv;�ۇ��R�I��x�s�j��P%���y��SO�r��xI�o�i�Uʻ_W�/���
PK�%���VJie�qj<q�����7e��[,�"��y+��v��	�fc�T2���tЗ#�X��'kgj3P��5�S�L�z���Pv�L��Ί4�EZ�5H���P����"�a������u��Xj�3Z�2�_��m^^���h�۲�g��nk�����T��z(:CeA[ԥ�-���e9��#)���.�*{Bk��:5��m� ���־�D6��SS��' $Ӽ��l�J�#��vng�k)��0A��}��1 h����n<EYi7587"<%��Z,�;��R��xJ;K#��W����^*��J���.>��[�����-w��K���>���4�˸n����?$*���/u~{�si���fH�!��0���n۵b-�=�
�<�����L7��^ �ʱb���߱�l	�W�pya��������+�
����`E6jU��.�֐S�R2�2!sƄl����1+ Ta�
�|�C����%����gO�6����v�2	8w�_Ki����/�gSΟL)����IR�s޵��V=<�T��'>����z[3CiBK�' �g�y�o�z��W�
 �ZѤbYf���=�����^�ƽ|��5?|�Wi̜H[�Z+��L�-;�tGTo�����E�u߄wJ�������rI�3Cs��I�LXTY]S��'��Ki��T�%����z,,`�jR�["�*-��GA��L{�`�-�z/�C�T�R��fPv�RR�uG�}k=�ѓ�Px�&�U�[U�U����Y��ki���R[b�K[�R�)�:/u��~��ݾ�P3�ք_���|Yr������?�z�g����4?q[�p!�ť�|K ��}�SH�ۨ8y����l5����5���?���x~���  �IK���eF���!��m/����y��Nz���г�������;�����<�xWP��@��Y󤏧X�+d�RL�XeW��Rk*��tD=^��%��i����������R���f7�Y�t���A�0N��st���6C��P<r�3�X�\� `��X���/�6ʀ���ƞ���P&Fd��N6��],���H��i�������N����������Oķ� ���G��w��~	iaҧ����.˿�d����&�TZ;B<N*�y7��f�M���G�X��+?Yŧƞ]�.�^A�!�⣴�͏Tتe��ײ�ի������z}�Wu����
h"̲`>��Dؗɫ��r�dNإ	S*&/��g�j�(�w8L�qQ.q�p�������S�Ň��ʴ�r�ʧ	��=�_�����WN��i*{-��|���~���r�0��	���	w��^�w�RI8=8�x\p}\���}������Z�ڽ{�ݿ�w�S��,���=,�	��D��,hMH�uB�ɋM�D�o\1e��.�rb�2A�k�+Q����c�i��~�wW�ֻ���-�N��d�x޷$i�95��Ě�sK��wAV��&a�=0�o�{�M�7\!�*)TD�6�(�q�nr�n�r�ׯ<���8����^�_k�
�gk��.tw�6P��2��O��/t~�{��S�[O���3�[���ew@��HE��}�F��7z������~�+XN�X���f`>bz�I��5˼�\�$e��I�i�z�b�E}7P���4�ҔT�����j|k�C�j}�&�,G���ꅔq<U\_/&*����4pݴ��6�c�F}*�����T� �#&��Z�u��Zunqs[|C
ٍK�Q�H�����5�m��
ǽ��vS!T�^�m�ZJ�۾�T.>���.��?�����C�,���#o�R�'�[�@���/�P2�_��SU����j�ai�;[��&kaZ���R����pk5�9Ϗ�$x.�+m?��O���#޾����6�ի�{�+|���k�W���Ҁ�r�um�>�S�������*6PD�]���p�i��~qUP+ �q��;�{�$��}Wn_�zpk��������y7}\���~��_�}��اtwH�����l��t���^���Ջ#ꬸ���)�N`͠�P�x��5�EЈQ�RFk%��u�_b�9����6L��z���X��^~���p��C���ⷿ�{s�U��g>j��`��p�O?�=}j��km~?D_$�}����\?�;�F�|��x�,f8���"g�����Ԅ�i�i^��+�
���r��;>&�%&y\=�]�pm{��u-�+�P�yʜ���M�Ȥ/{�ڏ�o�~��P8%3+��J�B����bG)#s��8�\v���)���xˋ|���?5���Η>�1(	��5�O?��?�aY�����I����iE�I[��XߢV�0�}h�o�ӽ���X#U" �/���i�-��ke�"�
WU������#��W��'�bC)���QR���(�$L����!>�b`�&ȑӄ[��ؕ���jŔn#c�D	�/���~�ٯ=y��������n�����ҧ_���$4��sϾѷ4��B?�a���{
����an3Z[px�����{���%Ǉ/��J��K��Z�k���bAkC&��^�M	�
�B8͋�N'@��i3/W�Zsx�����F%\�I���+���'�9#%B���d����)���pLލB��Z�l#Y}��	 2��4ٰ�4������k9��J�WA����>���8��-��7�������@�/|�ؽ�i\��h�G�y�����^�N��wf�ߩ�h�����Ui{�Z �Td��^��G��7mܫ��#��f���a�
}������J׆������,*�#� jC|��I��WhRQ�u�K���%d6�f���i���U����\���w��;O�}�c��̻>��/}�ݓ�s����p���7�6A ��_�E �VA�3�y��镯���t�.>Ȍ�6ײ���{ҖI*�r�2� ���s�>m�P���ٔ7��@��xS����]�>�
U�b5�UKIu�����e�i�GǞ�2��qA�x��y+RE`���{ΩW��(/�r?O��r��/Q��H��r��;���/E����=�;��O���`y������SO�vz[m�gAx*ߣ��Է�ջ"� �C2IUXUX��h��d5�㒮��R���Ůq4%+a����{�}�EM`B\���� �����MLPb7MP.>�E-4�4�\�����������������O��,������e���[Z��?��O �^�����>�j~��[o� <xG=]�u��
�>��{���і;m^��T8^�Z5u����54��mmV5�&�'o
�v�k�z#�����3!�U���(q#2��ܵ!o(��p�˔�g��I�.�,̩��2_'N��k����?���?���^�� ��}��F���t~��[��?�ҳ��P��׸x�S}����[h�Ro�N"����P}Z���[*8a�������խ����c_q��
���7�.?IB�,�m��*����>�0��וf�����m���5-˂��Jɨb�1S.Z�W%O��������px�s���/�{�ٷ�-�<�����o�� �g�ԧ���x�|��� rxn�,�����6�<S8�J�U��o"z��o�N�Ts���(��yO
�jz6O���"������
�6C����ܭ-nk�$))aۤ>�i�2"��2%%NB����J�f%>�
����K�ӗ�����qY꧙���F�^|I_��R�L�Uo{���ѷﷄfw�/|�v�j5��@� /����#K]�&�h�Y[M�IRQ6�g"�邈n�-�iOL;UL
ͤH`Ndc���X��J�d�G�*T�`�FB��5���B}�+��De�8-3��#�*�2�~�'�V�J�����<����������O������/�u�4��|��ѷ"�JT�}�8�M����p��~�N��p:ͻZka���:�D�ۙ���������nI�Q�h�k�y^��T91133)"�b��f��@�Y�Z�\r΀���W��X))1	@ں�-�1QQc�
�
�3���9�gN���U��N���,���>+���S�S^��N������¯��'�
�����w?�Y�؏��}�� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��1�Ӓ������   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X    IEND�B`�PK
     ���Zd��   �   /   images/a262aa33-74c4-460b-b0ad-c746896f6744.png�PNG

   IHDR   d   d   p�T   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  �IDATx��{y���u׹���Z�j��ez�����L�b'������2�eH$BaJ�@�dC��`�@��![G6NlϒqO{2��=��RU]{��ۿ�����1�'��n�u�{�[�=�s~�w��ʥ��1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�l�c@�a�z��Ti�R��)�|�H)����]ǧ0�Vg�¸K�F�Z���=:0��y��8L^a�&����4�"ϨH32ʐv4������>Y��6����=�n� ��w�H��)�~�����t�g��!�<T~V�Yz`�����j����ר�����Z�:@N�NF�ޢ���,S�ޠ��NY<�Zk��J��� m
& ̡T�nW���]����{}*f��>s���m�ݽ㯐[����u��)h~�����>�����R����h_�М�NݴC͠���ޘ�g>�?���g�~��P�R8葉ڤ+�T�O�8�,�`�UZ�	!�n�6�a���y6O"ǭVk��D o�D9~G��[�m���^�u�'^"�[^���O�N����+ DF�u
��v�����/M2�P���&���8\��
\��w�z��V�K3�K3���h㇟|������~ݟ����W���f�ȉCD�M"�!Y֕�.���n�Sf�	ch��G�&�q�H5���*o/��%�ݼIj��KI�Z����.J[�(�\ׇGk2�j�4���X:
A�tԿ�M?�Yg����K_����pkC通K�23�*0o�g3�$����0�v�g~�/+�W7��|��ּ�,un_����� I;���\��u��_},�~�n@"��-ob+b�v��X�I��f�L]�Һ^��U�8�E'?vV�x�C�k�;���M�}$�DLi�S����mQ�Ņ�:��(_Ug�����F�����	��ġ`VcrDqf*��q
4SU�NLm&U^�������G��i�8�3�.�۩.tؙ9|fp�[�D����W)�lSg}�����ѡ��0���%�]���pa�[���>PD���~󧢵�� �v���ԡ�����?�j�UZ��ε��@��_
��e���,�=McB�'�pt�&���.���
{^�K�zst���t��I��#���\N������r���4a�8&:��i�M����fS޻�0�*N�� ��%
V^��'B�%���w�1�@��Yuh$L�wQ&�0�3��	B8f��e�wA���Hi��%�?�p-,$|M^�0$ln���ÃN��'���S���;u���}���~g�| ��eP�>Gӧ>�����)3���I�+Q$d���򼴍�*ձ�aѣ�x�M�"D�ܤ,=E��Cdẝ��HKb�=~���kur��0!�-�)���!��D��)�px0D!�`����!��YҞ+sU9��x�T�J�,�OR@do6v�"�J��:������gB�K���E�����Ԡ?±��� ����s�Kh���+��7^mn����&]
wV�:{���i��u�Z�|�I��'��&��=�{��֠}m�r�<�r � ��c%ED��*�	���8k�0�Z��5�׃S�w����i@�g�ׅ�âz��w[�D'��I�Ar<��a�L*�އ\M����G�+�+��߰s[�����
��T�l1�z��=��.� �v+r�v��[�D�KO��c�	�K�N����[_|���S\�m#$ł��y��s��~)�oR�"�qm�ߵU�/�ԃpw��
"��U��2��Nڦ�<���w]B�^�X�U�F�ozZ�3d��(w�m����&�ҳɂ�d^J��)$��D� ]��X0�*\KIy,`Z�S�oا\G�څ��k�ԫ����G(4ED�+�i8���\r;Y_�Fa�bn���V�`���܉'�n��z �}G����#7��{�B���/ga�`:��v!{�%Z�A�q�P�w���~CYT�UM@u�C�D&�����m�O���KY`��Cs5�e@Q�f�\Z�m��-�%*$4�H`ٟ�i2WD�L]VCq�)�~�dQE�:�)IX˵喝
��O=E>U�)��:[[��Bβ�saȜF3�`H)E1��>>CN�?оs������=��;k�.�$�ҩ��x�~���p��_Α7�p�&q�@NTNu����	yф���ά�K���	]�WQ�6���p^S7����N�z��7e�WY��G�95�F��+�ÁBሚ�t�D�,UX�/��p $o�T(M{5�ր�2�gBrNa��r����
�7_׃s̟z���S��\!3X#߳�7��0��p�3��<��D4��Y���b4~�:��˝�7^�H,P��J�ܰ�K핛tv�y��'�w���y�����a2UNQ��8���/#z��!X�4Ee�w�.���9��� �ޙш���.U�5rI?��H�>��!���~�
S%6Y!
F��[ͪJ�亢�"PNтĚ�Ҿ��\�*Ȫ"�윬c�*#��%j��}���y�����﵌r+���Q����5��#w�<� o`Nٰ]M�꿞=��3������i#$�z,�Sm��}ݕ��}�{���ޑ(P���̄ZP^U<P��7�E�)s��p� �Jg�"L��s���8=�8�&Q&	�A@����d��U��Z%p@ e�w�C�� jT���xbn�[惟^��.�ӶxmhI�R�8��X[;��Dn�E~�^��WR# j.�5�RX�_�r�+��]�ʜ-��"���^�t늬դ^��G� x�s�⿸���ԉ?��Q���:�o��� j���g㝫���8��/�(���E�a���r��j�Tܻa/k8S�PY$����I:9s��;��1�M��0RE��<�Rھ��DR�y�2���D�*��$�ETdF�(�8*4�uD)1{6G�����@]-��=F���r��q����0��؜(y�s����@onm/;1�y�&�'����YH��.�KT]xP���SY2�A9qE���	r��������������έ����{>�����@S��/�c��eu��ʘ���	9%�Qڪ��x�"�4a�$ۡN�o��t���"��Z�m�O�ȉ�/SmΞ���%���b[�Ap�����29?gi�IH+�� p"��� xH_�\U�#�8 �=���� �Ʈ��Π�P|9�G�ex����)ݥT�$��5����)L��H��=�c-9Q��3�C���"��BS��4�=w9Z~j;�~����i�ě�}Ű"a��$�ڝ{<��X�1x;"g U.�*Y-���$�0��=��FG*��wi�f���zK�l^���~M��!t`����E�ޗ��5@���R�3�7(T�rl��<��T��;D5�PD��ѹ���d����\�p�!ё�I�#&��Hn=�Afa������[�M�����ox(�}��jߑ5*8�ҷ��D]�kduƵX���E��e��g���s5��w: +�KaS��q��0Y*rc�dZR��+J�*�G�Zc���"4A30��7���ޯ�Q�/�޸D���xs��D�p���.a����6�9%�3ա��XYn�"L[�˭"� �� 1��MR��(a�F��Pcs�6���w�UD#�ƴ�k�:&g�ɻ��P����]^[U��գ�W�s�%���@X���f�S�?��:	���.�B�r8�魐��57�ڛ'�G�͢�k�$�\.�Ӳ3�������|�R�|�|�܁�ڴ���P-���ץ�+Qhlo�)�^��˹!;�S��1C'�aT����Uz+�t�$½�;j�9�d(t��x����m�0H�Հ�"�Yi��BT������5���8R��/6�̽L�FKn�M_r;4��<�\�؊K�E~�%ut���ص;�2��e�@4�����*kY4S���X/���9������
�Y
p=���8�8,Xp��ͽʶ,�{F�>Q�H�Q�Ĩ�SCsnF���g���T���胁őX���}d�$PJR�_Ξ)�
���֠�hGh[���j����'M1��'�>�Hd�D5��8R��,
k"�Y!���C��\Ŕ�AqY�(7��=�b�H�Kr6���e�Nو+_2Kc�����]9ڪ�£���a�Y)@+[3N���?�u@Y�I��2�a^I
��a�|&R��e/Ki�Y����������<}8���$i��{{*2m��"��ZjF�R9\ c�YZ���V�#�j)y�*j�Pj�T))6�����Q�Ƥq��(؟���Z�K�כ�ό��bЃ�l%"w6�s9j�k^\	�m��J� ą�|�(�MҜ[_$9��.e�h5e��ؾ�eJ�F�M0>ߵ�����C���W��4n�&8A�{�^�U,|^x[]��~{�/ۓ��S���r�*��VM:�Ibh*,J2�{`PY��-s�&BU�S��!b%f6zx�"(���u��_NM��ϯ�]	p���[ِ�������C(A��ʚ�&V�%n��Ҳ��m��XZ)�77�lH>�~X���w>�ⴇ�P8Y��e�z��>�!,�S�}%�[��˕�P$+!g�0��Qd�F��-¬��X5�@�iPE�vٟa�T�r7����hޅme���-�a�����Ɣ��;GМ��`��?��{��~�ɿ��'�������C�r.r��Hf@�޾�ѹ���J�ƲЛ�J8����1��� B.N0���=6ۈ3ei��0����E+<÷�V�sI���ϋ{=)�[Q�����#�Ap$�r��q�a(�`�FQО�Y��jî1��X�~�ʍ����C��V!��e���z�3�r�[)W�`�'��?�%��_x���gg�~�Gk�7l>�UH��E�ǡ.J!�dv��:�Ք&�6N���&�1�Ri3צ��=#*�!>�
�mI��P�{�0$j����쵲�ABf�Y֒#����j�����K+GDA�iy_dv�Q��M��T�b���xm.��P�vű|����g�e�X:�JP�W�})B����qQ���H��=���t{��?;�U2�1�	���`���'�~?l.���!Q�w+gD��w��<F��8� ��#$�I�G^�Aa)�un��-O!
c�	����ԋ
�	i(6;��R��	�����|#M�RJd�sRa��
VO^'ANL��Y�k���PY��6��Z��<mMf7�4�t&{,E)�*v�t$F[��1!,�Y�y�s������}2;7YW�����c�q�u�x��T_,.y�}?}�y��,�Ӱc���Z��团�`����)&��|,Q�%�3�Z�T���OD�R����M�όy����|DJ�s�<���O(]��Yx�L�|��X�ǀ�ANY�ؘ 2��H0/n]��z�̍�s�B$+D���"Ys3�T�
Z9?�`NY�h$�(ͲQj�cIQe�_�)��T�~.�t�̳�z�U:�����!�����(��+/�����_s���n�E}��P�{o�����\P���r���J*@S)GG����Ae!ȋ�G\^���P4l�ݞO��+�;�,�}!<��F�R�L���=T`��v������[C�����8/QV�I��@�[�%���-s"� d����uH2��<�P1��:h��gI>�b��I�ѯ�Ch5�������7���st�]��\�v�~7-_x�K��c����YtH��O�-��:�F�"iK�\Ŀ�׏���4�ϐ�x��
�d���Y���Oi+���V���!���h�w�e
 Ң)�;�YِR;@nom��@O���#&���V��UBq���ͯE�.E��4�΂+�5YO�{�F��`d�mp_>��A�Q/���t���h�(��;�_�Ï�|���|����k����W�n�u�1��H꿡������H1��;�^�[��dQ!G��Ȇ2�@qN��A!)�k�ҶVE�V��u2��f�u�k$xn��(0p��]6�F�DSFF!^���+
��l��?W�yn��\Ԡ)v(�6�r�u$��k�
PEO!���$c��'�,]
�Q=�st�t�\���ׇ^�������yo����G����!�v@fg��k/����?���������S�ҡbЅ��e�~i+e%BVG��b�f�n��Cb,�N�w���Ƚ �T�k\�K��'���V��h���]�B�� ^�>]�����lM+�wJ�2u������5)Ly�2�MR�UI5�}��L��k1����k�	oN9Vy�߇�#Y1a;T�&�.����í�~��c������c��i���?0��e|�)�u�T���[itď��FC��'�Oūx��i�\�s����3Μ�-���'���*��jו�6$���-��4��"k����z��J�Z��sը�Pvo]B5��\Q�{߳5�[%g��ٽ)8�eC��0�,~F�_�J��@t�4U�*(�R��#��>�M-�hQ�3�܀�t�m�e�l�a=^s��������~�wx�̇�w�������K��|�vV.��}�?���?b��;����"�e��=�f/.��kT_���En��u:��!j֏H����V��|W;^�K���MD���*��4���AUy���Ss)�f������|��#;���.�u ɎHw���.!��#К��BZG�����8�%��N5O�zGSY�u'�}����O\B� ��Ȯ�H�N���a�'.j�.Ҝ�g)�#p+Ti-Qe��E����a{c��n.�������ճF��w6�S'�������:���H�}R�sn)���>���z�&�3�Uϣ�?M3�����Go�V�3����W_s+��&��N/�G�+���Q���Yz���k۝f�f�����@{��㙄�"����Ju��9�r�i�v������������X��� �:��LT��N{�/)<L����l߭;�f�y�5����ߗ{�<r����.��y/��^"�@�ZI=�F?s �<8^0��U�s���t�s;���H�}oJ��y�V_y�q�����d�����~�v>��n�%G GS+]A1��4��x*�������D�ۊW�=W��k�>��/]�򯷛G���	��P�_'�*�.kqgv{��RoQ7�d�*qR
}EQ��0�і���|�>9Bൕ�e2�-�i��,�bؕ=>'K�w6h8�KG��� `<PRvP<�)���y���?�ɠw��G%�:��=SSt�0Eu�婙�H�Z��S�z��M�yם��?[�N����s�<E5�X�����w3���}ȁG�CwΝ�J����is��*4������V��6}���ȼ���T+�����ڌ)	w�9�_����W~��W.�C��%ZlP-h������}/^�L?N/|�b`|P��֚l�nܜ��U�y�ؗ��ڇ2�[��}�[����<t9`@K���w:�W_���BՇ�{典H�o�4�f��2-��_���[�p�C��
��9.'u!\1���tz�5|�|��>t���W�9��D<����Auߙ'�~�s�"�?�7i��D�����G~��_{)�]D�D��.
ɵΦ��j[Mz��ץg�͆t����q����r�N<�m�W.~���CTi�݋�%�W�ƉluKu�P����FS��5����� ~i�~��wt�?�}�w�����O��O���wf��c�W�c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2f�D�{��w��    IEND�B`�PK
     ���Z"1^FHo Ho /   images/4efcf596-32b1-4e3b-9735-2bd5fa764fde.png�PNG

   IHDR  �  �   �r��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ��IDATx���1mA  ���+w!`0�t ^z )�-(R^$E�}i��_]���s� ����\k�       ����|��5 ����cp{��朏��s p'         �%�          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��     ���<F��~��k�fq�\��PVeqU������T��T��aIl���6�4���%��5�j)mm<j�j����J�"" �s>�V��@X�3�x$��?;3���_�y}     � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	���7�o�=���������r�l��ʲ����1(5���z��7       �Z�vm�1�@����}����c�3?�7�۲7�S���?p��͹.x�%K�
���q�GF]]]6={��#�8"�u����o����///�~>�y�>/         ��k��o��F�ڵ+���Ν;���cǎؾ}{6���Jl۶-{=I�~s
^E UEEE444dӫW�l���ߺ���UUU         t���ټ�bڏbϞ=Y�e˖x�嗳s�l޼9���g�>�;�\.�썍�q��G�QG}����޽{g�         ţ�����z�󝝝�u��,tߴi�[�q���}���������������c�9歨�v         `��r�^�ze3x��w<�w��x���^Ȃ��lذ!����ަ��>�?��8�㲨=���#          TEEE{�ټݫ���ׯ�b��������6x(UwJVuuu������          ]�{����ܜ�~�v��>�~��l�}��رcG@��S2�8�,b�O���������          HEMMM455e3al���/�O>�d<��Sٹm۶�b%p�h����'?��2dH�766F.�         �B�o�d~�<���M�6e��ڵkc͚5��+��;E#�����YО�UG>j///         �bҧO�lƌ���y��,t_�jUv�ٳ'�P	�)huuu1t��lN<���          ����!��ڲ��������}��ձe˖�B"p�����/ZZZ���'>��z         ����ʷ��mذ!���X�n]tvv�L�NAhll��O?=N;��         �ֿ�l&M��ms��b�ʕ��3ψ�I���d����)���E�MMM         ���իW�;6��_~9�ꞏݟ~��T�IJ�޽���5���\.          8�����7o�U�V�_��X�~}��$p��ѣG�1"�          �NCC�[����?+V��Gy$��]M��a���>dȐhkk�SN9%���         �ë_�~�L�:5֮]˖-��<�����t�#�<2F�g�qF�m          ғ_f��ܜ���۳����}�ƍ����C����[[[���,          (=z�c�f�nݺ,t�Gb������C�gϞ1r��8��3���>          (l�|6ӧO��+WƟ���x���;�	'��ƍ�aÆe��         (.�����֖�ڵk��{�������q�9(�!�СC��sύ���          �42$�M�6e�z�سgO����TWWǈ#���}��          JS�>}b�̙1q��x���O�S������RWW���q�YgE���          ���)S����_��{^z)�����Y�����ڢ��2          �TWWg��?��X�zu�}�������;Jccc�{�1r����r          F�=mii��g����+�zꩀ�"p�}����ĉc̘1QVV          p�����_�B�Y�&�׭[�vw�S�޽cҤI�v          ����2dH�^�:~���Ɔ��C�^�b���q�gDE��          �F.�����:th��o�%K��K/��63����7n\�;6*++          �B>t?����SO�B����7�iӦ�4	�K\MMML�81۫��          �����a�b���t��رcGPZ�%*�`�ȑ1cƌ�ѣG          @
***���=F������{��A�^�\pA80           E���1}��3fL��W��U�V�O�^Bz��ӦM�6��7�         @����W_}u�Y�&n���ظqcP��%���2Ǝ�'O����          �B����_}<����t��عsgP|�E���%f͚���          ����<[�<r�����<�@�۷/(�"�����͋N8!          ��t��=fΜ�G������nݺ�8܋L�[)�sNL�:5**��          �����c���q�w�믿6t���^x��	          � ��E[[[477��ŋ�'�
���TUUŔ)SbܸqQVV          Pj��k���+W�/~�رcGPx�N��s�F}}}          @�;��bРA��_�:~�ᠰ�TmmmL�>=��          �_=z�/�8N?��X�xqlٲ%(�4|�������.          ��6t����W�w�yg,[�,:;;��	�HMMM̞=;F�          ��֭[̝;7Z[[cѢE�m۶ ]�1p��X�`Au�Q          |4'�xb|�+_�[o�5V�Z�I�������<yrL�4)�          L]]]\u�U�|�����c���AZ�	�������hjj
          ����r���'�pB��'?�6��'jԨQ1{�쨩�	          ��jll�뮻.�.]��sOtvv���=1ݺu�9s�Ĉ#          8t*++c�������-��[����=!������իW           ]#�_���ӟ�4�x����'���-f͚�          �juuuq�5��=��w�uWtvv]OM}��ok0gΜ�ԧ>          ����b	�����rK�ܹ3�Z�èw��q�W���          @ZZZb�q��7�ƍ��#p?LN>��������           �ҧO�����zk�X�"��.��m����cڴi�5          �������KcȐ!��_�2�x����w�����袋���5          �����G}t���?��۷��������/����V          @a4hP,\�0~��ĺu�CC��������/�nݺ          P�z��_��cѢE�bŊ���bcƌ��s�Fyyy           ����2.��hll��K������r1eʔl          �Ɀ����;�#����C���".���1bD           �i�رQ__?��c�����'p?Ⱥw�W^ye4(          ��6lذ���?7�tSl߾=�x�QCCC\s�5ѷo�           JÀ�뮋�}�{��/N�~�80��ꪨ��          ���e�K_��o�9�|���������������           JSmmm\{�hѢx��G��N��1><,Xeee          �����lyvuuu,_�<�h�C[[[̝;7r�\           ����y��EMMM�w�}��'p?@���1k�,q;          �.�������"����w��#p? &L��ӧ          ��9�󢪪*�����	�?��lʔ)          �a�lWWW�m�������&p����"���          �����=���c���"��!p����b޼y1f̘           8mmmQSS��rK�����	�?@>n����O?=           >��ÇGEEE��G?�������r��vq;          p�����%�\�E�����K��?���ٳgǘ1c          �`:��Sc�����,:;;��#p��M�g�yf           
�G��]�v�m�����{�:ujL�0!           ���:+^{�X�dI p���>;&O�           ]aҤI�{����	�ߦ��=fΜ           ]鳟�l�ݻ7���(e��o���1k֬           8f̘�v�e˖E������5�ϟ�\.           �|�<w��,r��G��|�����^zi���          �ᔏ�/���رcG�Y�&JMI�q�e�Eyyy           � �7_q��o|#�{�(%%�y���}.jkk           %555Y����=�l���$�����ꪫ���>           RԳgϬ{��7����z��������K.�          @ʎ;��⦛n�}��E�+��}�̙1lذ           ('�|r̞=;/^Ů������Yg�           ��3Έ_|1���(f%����Ĵi�          �������'{�(V%�80.��(++          �B���b���o}+���E1*���G�q��Geee           ���������o��[�F�)�����<��޳g�           (�%��N����v�ݻ7�IQ�3gΌA�          @1ijj�iӦ�w�Ťh��#GF{{{           �s�9'6l�?�p��܏=�ؘ7o^           �9s�����c�ƍQ�.p����+��2���          ��UWWg��׾��عsg��
�s�\tttDCCC           ��>}���_�������3
YQ���g��O          �R���'N�?��QȊ&p6lX�{�          P��N��ׯ�����Q��"p����V��r�           (E��z��q�7�֭[�|��.���֭[           ���ݻg}�w�����BS����ɓc���          @Dsss�}��q�}�E�)��}��1iҤ           ࿦M����?cÆQH
6p�������(//           ����"�o���سgO���gϞ}��	           ޭ��1f̘��v[���O=��=zt           𿵷��O<�V��BPp�{�^�b޼y          ����r1����b��푺�
��܋.�(�w�           |��������w�������
�'L�C�	           >��N:)������L�޷oߘ2eJ           ��M�>=V�^�7o�TD����b���QYY     ��ػ�(��;��)00�.��4�R#�A��c�&z�9ɉ���$'�����I�;!ш�b7�=XŀH�D�I�����DQʔ;3��9Ϲ�/1̝�e���     _ݺu��+��o�1�����Z�i~׮]          �#WRR���_=rQ��M�6���??           8z�]vY̙3'6o��&��+��"�ׯ           ��%�\����"��t��F����7           (?C����z+f͚�$g��+��K/           ���_|�A���F����=��5
           �_������Ϗ|0rEN�%%%��{           *�i��3f̈�F.ȹ����(������           *N궿�������سgOU�qr/p?묳�E�          @�;��c��SO��S�V�%��f͚�g�           T�s�=7�x�زeK��9r*p��⋣nݺ          @�)..�"��￿J�9�w��%           T�#F�K/�+W���?CN�yyyq�e�e�           T�������K㷿�m��r"p6lXt��1           �:%%%ѷo�x��w����<p�W�^�w�y          @ջ�Kb��ٱ{��J��*�ǌM�4	           �^�V���N�g�}���J�}��          �i�����cӦM�z�U������U>D          �O�W�^�w�yq��V��VY]ޥK��۷o           �{��?�|�^��������??           �M���1f̘7n\��g��%%%q�	'           �k������OǊ+*���$p?�s          �ܖ�����w�qG��_��{��nݺ           ��_�~ѩS�X�dI��W����}           ��ԁ�3&n��
��J����           T}��Ν;ǢE�*�~*-p7�          ��:��s㦛n������}���Ѿ}�           ��9���{��1o޼
��J	����Mo          ���?������+��WJ�>x��8�c          ��k׮q�	'�|P!_�R�Q�F           ���ѣ�o�޳g�h߾}           P����+k�W�XQ�_��w��          j��O?=&L�P�_�B�T嗔�           5�����G��?��\�n��G�����           ��(,,��#Gf�{�~ݨ M�6�           5ϩ��O=�T�����׬�����OϪ|           j����6lXL�:�ܾf����ՋSN9%           ���8�x�����\�^��#F�����           5W�-���1cƌr�z���ȑ#          ��o��ѹ����y��          @�שS��ܹs,Z�訿V�rJ           P{��<���-[�	'�           ����z(�m�vT_�\�#FD^^^           P{ԩS'/���Q}�r����c�С          @�3|���	����M�4	           j��;F�bٲeG�5�-p?�S          ��+Mq�ӟ�tğ_.�{��ͣ��$           ���&M����#��r	�������           ���_�~0 ^{�#����S�~��'           >���޽{GӦM           �t��ڵ�U�V��u�>lذ           �}N>��x����*p/..��={           �3p���4iR�ݻ��>��~��Ea�Q�          �i֬Yt��9.\xX�wTuz��          ���޼���FIII           �?K��C=eee��9G����?


           �Y�ƍ�k׮1o޼C��#�SM           3`����5jݻw           8��?��QVVvHD�{�����           ���7\}�ܹ���G�80           �������&M�D׮]           �H�������={�|��v�>`�����           �"6�����={�~�a����           8T�{�.���~��ѵk�           �C���'~��V�ޫW�(((           8T-[��֭[ǚ5k>��+pO�<           ��={�_�����Mp���m۶^߾}{�ݻ�S�N)**��z�YV�^�          *_�ѧM���sȁ{�Ν�A� Gc׮]�iӦ���c��ͱe˖غuk��p}�J����Ǝ;b��ݱs����={����N�:�J�{��������ׯ���o�{�q��ѨQ������u 
         �w��{�%<�C.�N<�� �ϓ��6dk�����/jO�zUK?���I��*E�M�4ɂ�f͚E��ͳ۴Z�h�ݦ8         �?u�֍nݺŜ9s�1w K��?����裏b͚5ܦi���)�W�>��4l�0Z�j�[�>���c��y         ��z��u�{
�:v� �7n��U�Vp{�S�k�-[�dk��şz_��޶m�l�k�n�m�         j��={~��)p/))���� �fJ1��e�b�ҥ��%KbӦMA�HS�Ӛ;w�oO�{�P֡C���{Zyyy       �^�v������ۣ��4{yϞ=��;w�ݻwǎ;����y��ԩ��}�ի�@�����������կ_?�ur= G�c���-[�ڵk?�������# �RX�����hѢ,hO7T���ͬY���O�F��S�Nq����_�       �����6d���͛��~��[�f�z��sɾ�=ui5l�0�6m��6n�8{9�k޼yR�@-�����⋟�>�;@VVV+V�����g1{Z�ׯ��t���{�e+I�����w��%�u�mڴ	        ���}͚5��裏�f#��7fa{��^]�&�ɻ����f͚e�{�-�պu�hժU�� ��Q��J�!@�KA����c���p�;wn����c�޽�z��l���k��҅`��޵k�())�:d!<       P�R�����=[+W��?�0��S�^ZZ�#�Ok�ҥ�z_�Ҕ��(��]�vѶm�l�	� �\�wK?R�Ͼ0p�޽{ ��V�Z��~̙3'�����I��f��V���J�{:���O�vA       G'M+_�lY6|0�i������5�[�.[i��'g�{��۷o��;��c���( ��4h�=Ƨb�L�P�lٲ%fϞ�E�i�c���6o�o��f��6m�d�{Z)|�[�n        �-E�i��%K��im۶-�<����O~~~�Aw�q�J'�w��Q�PMu��M�P]�ݾ��n���{1o޼سgO��Jǟ�5mڴ�S�Nv�K�޽����1_       P��ر#V�X���,�ŋg���=iZ��ի���odo����=MyO]D���� r[
�_x�O��s�F�E�֭�ʕ����}�̙YԞ�a��k׮���|����}�{��      ��n�ƍ1���+��ij;��'���ӧgo+..�B�N������[� ��!�n����b�����E�bƌ��[oŦM�*Zځ��SO=�Ms�ׯ_0 �t��9        5Bj0� �>� �׬Y�l۶m�Y�fe+)**�Z��D���C��#7n�Z������܏?�� ���޽;fϞ�E��	���������c�ԩ�jڴi�4H�      @��N7_�`A�ϝ;7�-[fB{-WZZs���֣�>��;w�b�����T��x|X�{� �W�`Z�pa���曱y��\��c{��լY��߿6�=�       �&�qi��{ｗ��i� L
������-[F�^��O�>ѽ{��S�N P9�@��ӧ��ѡC� �|�Z�*��׿fQ������u�d�c�=6C���w       �
eee�|���Q�ҥK��ڵk�Lq{ ػw�l`ӦM���Y���o�>�֭ ��۷�[o����ij;Tw+W��?�����#�dGt:4N:�$�       �p�v�9s��̙3��wߍm۶����l�t��z(�,�N�O}D��@�J�zQQQv��>�Ӄ2 �o�޽���^{-�y��I/�4������dS�O>���رc       @y�Ϙ1#�0v��PYR�hѢlM�4)ڶm�Mu8p`�2 G/???:t���������5�Óv�I�S�N͎-��"���wLWz�p�)�d�{�U       ����,>����>}z6���]�*�^�:��l�݇�Z�
 �\�N�-pO%< _l�ҥ���/gU��Sۥ~��4hP�92�=��       �ϓ&e/\�0����o��͛r�'c�4pȐ!Y+Ѹq� ��w�q����{aa��3 >G
�S�>mڴX�re JG¥�iu��=N;��۷ov�       �f͚��_���6TG�N�4)z��'�|r���'


�/�σ�?3po߾�V�ϰiӦx���^�-[����͛���-[ƈ#b���ѠA�       �vJ�g͚�M�;wn6�j�={�d��*..�ĩ������ �M�6Q�n�عsg��g�L�dɒ��_�o��v�D8|k׮�ɓ'ǓO>��TNS�[�j       ���H�g̘���5ٶm۲Miu��18dȐ(**
 ����{l,^�8{�3��P[-X� �y�lW%P>v��S�N�iӦE�޽c̘1ѩS�       ���7���矏��FK�.�֤I�bРA��|������{*�j�t��{�O<�D�s��{m߱\]�t���:+���       T�W�Φ�O�>=�o��?���Z��0 
��k߾���?�Q�m۶P��޽;^{�lb�ڵk�<i��m�ݖMr��W�}������       ��H���Ν��Ꝇ�ׁϖZ��z�8����N��M�@m��~�S�{z�,..��"��o��VL�2E�U,��0v��h׮]�y�1d��;      @�+--�7�x#���lr;p�6oޜ�L�?i �Q������&5c�~�;j������'�x"6l�@�X�jU�?>��K�����#???       ��q���˱m۶ �\j�f̘���ݻg�DϞ=j��F�F���?w��ٳgO���Yؾq�� r׾���瞋��;/۩      @�Z�v���}׮]��y��e��c��ѣG��c���>��m�6 j��{���o��<�H�Y�&��cŊq��gGp]p�QRR       T����4��7ވ��� *�ʕ+����=�X�~��q�)�Dݺu��J�g�mڴ	�����ߏI�&������/^���o�G�q�Fǎ      ���hѢxꩧ�����kݺu���f߇��zj�5*�ի 5�1���
܁-Ű?�p,X� ��#mZ�;wn0 �[�l       ��}a��Y��z�7o��<^x���,tj�V�Ze��EEEѨQ� ��6l�O<�D���+vC����z뭘9sf�;��sύ���       ��,\�0�L��rϖ-[����_�"������kݺuv[��o����ꪴ�4�}��x�gb׮]�|{�쉩S��믿g�yf�~��QXX       �U�Ve��3�}i���ɓ�^j���q�i�E�:u��jٲe������PݤI�/��r<��c�7��ٺukv��ꫯƥ�^�z�
       �غu�⩧��~�ZVV@��&��f�^���>;��� �Mz�j޼��'�T7K�.��'ƢE���?�[n�%����]vY��      �O۸qc<��Y؞N������ǽ��S�N�.� ��� �M���`@u��5�c��M��Mp��Y�fŜ9sbĈ�E[QQQ       �s�ά�x��'cǎ�,�V���o�=:w�_|qt��% ��Գ���� �.��.��L�۷o��ٽ{w�+��wމK/�4���       �U ���oǤI�bݺu�l�-�믿>N:餸袋A��Գ܁je����1:K�,	�C����;�O�>�}-Z�h       ��ܹs㡇�+VP{��-3f̈Y�f�g�g�uVԫW/ rէ�f͚@.JGc=�����s�e��D�XK�h3z��8�쳣��        j�6�#�<ӧO��ڵkW<��S��k�e�܇yyy�kRϾ?p/..�+�I��NL�81��8Z�6̼���o|#:u�       5��ݻ��_�G}4JKK ���c���1mڴ����u@�9`�{ӦM �l޼9~�a;��
�|����/Ç�K.�$���      �&H�[?���v�� �,K�,ɺ�4���/�F�@.HM���=�s�3f̈��?��*�޽{��_��s��UW]ݻw      ��j�ƍ1q�Ę9sf |��M��iS�E]�	�����TXX��{�&M��mڴ)��~�� �,}�Q�����i�      @�TVVӦM�G}4JKK�pl۶-���x�����_�z�m�6 ������@UKS���غuk T�}��?�����ꫣs��      ��-[���K�.��1����Og�qF�{�Q�N� �
��ƍ@UرcG<���YX
P�֬Y�_}�5*�?��(((      �\�&�����^x!�P����<�L���;q�UWE׮]��	܁*�dɒ��{�� W�����ڼy��k��֭[      @�HS����?�-�
���o~�>|x\r�%QTT �E�T��>��s�裏f�� r��ŋ��?�y\|��q�)�      @UڱcG�ZL�6��v�¥Ǚ�_~9�̙�Ms/))	�ʰ?poذa T�u�������� �.�ѽ����~|�߈���       �l�g��~w�~�� �L�������iH�i�@E��7h�  *ڌ3���m۶@u���D�k��&�u�       �a׮]1eʔx��gMm�Lz�y饗��6��ַ�K�.PQ�)M@����c���P]�I7�pC�92��կFaaa       T�իWǸq�bŊ��4����7q��gǘ1c"??? �[Ve�׭[7 *¢E��������K;��N��=�}�;߉-Z      @yJ��|�W����;w@.)++��<�̙�\sM�j�* �S�7k֬(/// ���/�'N�ݻw@M�dɒ�����ճg�       (�7o�	&�{� �,���~�_~y:4 �K�7mڴ^ ��]�v�������j �T[�n�[n�%F�^xa�0      �ٳg����شiS T;v����ǬY����F�����@9ٰaC�q��tc��.��3���ի�ꫯv�      �4Hp���1mڴ�w� �͌3b���q�5�D�n��hd�{qqq� (��͋��+;.�6I;�����;����h׮]       ��+W�=�ܓ�Tg�ׯ�n�!F�_��W���0 �D��QTT$p�J�=����#�<eeeP�Y�&~��_�UW]      �����/�ĉc���P��l�ԩ�lٲ��w�M�4	��%p�ڎ;b	���o@mWZZw�}w̝;7.���(((      �OڵkW����+P-X� ~�ӟƷ���8��p�ܝ�?�0Ǝ�W�j����hذa�۲iӦ�z��W�ݘP��I��߳�ȍ7      �dÆq�wĒ%K�&ۼys�x�q�ęg� �*��֭k�;p�f͚�ƍ˦S}իW/5j4H�X���!�ԩ��~�����y��׏���O}Ϳ��o�q�ƀ�n����_�"��_�5�;�       j�y���]wݕE� �AYYYL�<9V�XW^ye�|�;pD�d�?��O�rS~~�����mڴ��m�F˖-�U�VѢE�,lO�zyK�!p�H�������k�_�~      �>��g�}6y��P+����jժ��w���K �'��������<[��w��%N<���ڵk���ѡC��رc6q����}���C:�"18f̘8��s      �=v��&L���~; j�4��g?�Y\}�Ն�k_�� _`׮]����>�z� w����N�=zD�n�8�gԨQU�gJ�;p�}��D�+��"
      ��>���;vl�^�:�Q�F�Ջ�?�8��J�~Ґ�ѣGǅ^yy�U�Ӳ�����#�6o���v[,^�8�z��q�}���^�zEQQQ��;\:Yaݺuّ[���      �fJ�� �t�35Gf��֫Wo�˩�(((�n�`�t[\\4�VӦM�y����������?P��!��<�L���k��O ���yyy�pk֬�[n�%��j�m�v�ްa��Uw�|s�΍_���q�u�E�f�      �Y���x衇����!��-Z��V��4i���"���p=M`?�
�?�f͊_���o��oѦM� �'�����	��gZ�pa�~��e˖�j���={������:Hxig�����l�V��_����}/ڷo      @�WVV'N�_|1�=�e8��G�1��شiSt��)[�s�Q��"�yyy6?�������W���~��ѽ{� HLpꭷ�ʎ�ڵkWP�:v�'�tR�x��qV�M�q�|�� n�ƍq�7ĵ�^�"      ����Ҹ�����rG�WRR�E�)d/((�ޞB����4>�����[��M7�W^ye:4 ���IO=�T<��v�V�t�U��~��'W�cw�ph�m�7�|s|�[ߊ���      P�lذ!n���X�bEP�RD������7�t�?j�i����{��l�~�w��j�� �'S�L��<�<͚5�dۋ���&H�;ph�Iw�uW\u�U�/})      ��c�ʕq�-�d�;U'???�v��{��&���=W��b�(c}��'cݺuYC������~`��ᡇ��>��۷�aÆeV5mס�OYYYL�0!v��#G�       �͙3'�����|T�&M�dQ��A����M|��_=>�����w��������V�{��ꫯ+���|:4;��r1�/m4z���c�F�      @�z�W���˚*W��|�	'Ā���lѢE �o�ܹ��_�:���h֬Y ����?5x���A�IGa��ib{�֭��KO,

bϞ=��?��ñy��袋      �-�wz�'O�g�}6�\�5ʢ���GqqqTW�¡Y�jU\��Y�~�1�P{ܡ�KS�Ǎ3g�*F�%|�'�i��V�vঠ�y����Gp��y����/�v�      ��JC���?�k��T�v��Ő!C����G��7nEEEQZZ��[�n]��W�����N�:P;ܡ۹sg�;6�̙��4��W�^1bĈ��GK��w8r)r߾}{\q�"w      �bi���~���1cFP�Rw���/}�KѦM��iRK��S_l۶mq�7������ҥK 5��j�����o��s��+E��k�ȑѬY���Z�j��~ G^�����oֈI      P�����w�y'�Xi�y������I�&QS���w8ti@�M7��^{m���#��M��P��v�-�ĢE���չs�5jT�m�6�Z;���믿;v��|�;QX��      T�4�j�ر�U���СCc���Q�^���R���x|뭷Ʒ����ׯ_ 5�B
j�H��Z�.]������g��:u
�O����w�}7ƍ�E�&�     @�H�����A�ٴ�!C�D�:u��04�L:Q㮻�o}�[1`�� j&�;�";w��v����O�ƍ���O�>}�D^^^p�t1����ݻ7��7s�̘0aB|����      l۶mq�M7Œ%K��W[��}Lp�#�gϞlH`�:lذ j�;�i��w�����^��JX#F���u�����(5j�6m
�|L�>=


��+��     @I����c�ʕA�*..�SN9%���7_KC���eee�����?�1��ӀR�f����I;���Θ={vptRLڻw�8�3���|���X����W_�z��ť�^      @�Z�~}�����5k��'<xp><�}gm���&M�Ć82{��|0�o��sN 5��j��Sm���1k֬�褝�g�}vt��%8t)p_�hQ �����&�@     ��v�ڸ��ȝ�N�0`@�1"6l���T���M�2%��P@�!p�,�P�����7��\�:ubذa���|4֑Jc@�Hh�1��3�      ��lܸ1��.n/?�;w���:+Z�n|Zj*�ϟ��KEj��cP�)5�{���W^	�\III|�+_Ɏ���ܡb���Ύ�;��S      82�7o�o�1����K�@�խ[���Z�h@�IE���8� �7�;�P�'O����/��iРA�=:����;T�tZ���ߟ]���&      �óm۶���c����ѩ_�~�92������T@�KCaӠ��ÇP}	ܡz����g�	�LϞ=����"w�^�F����(JKK�)r���{���E      ��ٱcG�t�M�lٲ�����E�>}�a�z�C'p�����/k(@�$p��W^�)S���q��q�9�D��݃�.b��ʕ+�8eee���.6l%%%      |�]�v�m��K�,	�\�6mb̘1ѡC�����I�i�P~RC1~��,rO�o��G�5��ٳ��g�4�=]l�O��cϞ=q�wď~��h׮]       �m�������͛��u��ȑ#cȐ!�����T�X�"���;�3��_�%kÀ�E�5ĪU�����v�q��.�Q�Fŀ��ӢE� *���۳)?�񏳓)      ��;�o�[pd:v��w�����w��63]w�uѭ[� ��;� 7n��o�9�9t�;w�.�@ Z	�nc��]�6n�����~��      ��޽{c���1cƌ���$x�I'E^^^p�4P�v�ܙ5������9@� p�jnǎ��6�&�5bĈ8��S]lUcP��.]�ƍ�k���q�      ���w�}��o����$ƌ�5
ʏ�*^j�� ����Ѷm� r����td�=��˗/M�&M��/��;.�<�8�ئ��@�5kVL�<9{�     ����'���_~98<���ѣGǀ��'p�ʱe˖��[�'?�I4n�8��&p�j���EM�=��΋������� �5k�֭�r=��s�&��#G      �Vo��V<��c��I/���h޼yP1�[C�r�v��[o����� w	ܡ�z���^�X���:�4hPPuҎc�;T�|0�G��}�      �6��Ϗ����޽{�CSXX_��cذa���T�Ե4m�4֯_@�[�ti�7.����ls	���P͘1#y�����d.��lG1U+�|�A �/��Ogir�N�      j��>�(���ؽ{wphZ�j_|q�i�&����C�5kVL�4)�ʀ�$p�jf���v��;fOB6lT�t1T��;w�رc�?��?���      P�mݺ5n���ؼysphҩ�cƌ��u��'5�������/ɾ�F�@��C5�.�Ү�]�v���:�����Ow�L�C�۸qc�v�m��(�ԩ      PS��"�nl͚5�KA�9�}��	*���ƃ>͛7�6� �E��DYYY�u�]�aÆ��
��s���#�#̀��lٲ���{�ꫯ      �������b��kӦM\z�ѢE��jܡj�&oܸq���?�?�� r����I�&9��4j�(.��h߾}�{�ի6�-[�P��O��:ur�      5��ɓ�7��X�޽�A�i�;U���:;wc�Ə�cߋ�C�P̜93������9昸��ˣI�&A�J;���1[�ڵ�N8!      ��x饗��g�>_~~~�v�i1|���5h� ���c۶mT��?�8n����я~�����	�!ǭZ�*Ə���g�ѣG\t�EQ�N� ���}ɒ%T�t���w���_�͚5      ��.\'N>_�F��K.�:�#M��C�I��]w������M@@��C۱cG�C���4�lC��3�<3������-�7o�;�3~��Fa���      T_i�n��מ={��k۶m|�k_�&M��%\�|y UgΜ9��c��\@�R2A�J������ի�OKA�駟j�U�V�ŋ��ɓ��K/      ��RԞ�ȝ��ٳgm֩S'�=�Bnx�駣}��1p�� ���r�SO=3g�>-MN\�z�
�����=�?�|t��%      P�L�81,X|�4Dpذa� ��2�IS�a�`�֭[G��w�A��~L�2%��z���W\��C5��8K;�w��@n�0aB�k�.;�      ���^{-^z�೥��_t�EѣG� �	�!w����;������P��c6n�w�}w���JO����8�c��)�OGj��� ����Ƹq��'?��#	     �V�X���ي���k_��!��D�f͢�� ���@�[�vm��]w�u���@��CIǛ�?>�n�(M��ꪫ�8��-�8�CnJ� 8iҤ��       ���b�ر�s���Ӛ7o_���u�H��S䞢Z 7�������O��g�@��Cy��b�ܹ��R�&��ȝ�ϑZ�ۦM�%%%ѯ_�      �\��s�=B��h߾}\~��ѠA��zIM��א[{��ԩS�x�T�;��˗ǣ�>�M�6��v]5��r߄	�c
�T      �5���={��c�>��:�Ï_��Җ����e�K�jX�l��j�؊�=��˼�8�E�v��$��E�U�UHt$$!�*zG4�����h�([���g�_$v{�9�>�뺃ˍ3&����:����򣩀ғ��~��_����0`@ �C�%���1~��_GSSS�aÆeq{�޽��p��w����p����,*++      J����c�����&L��=�XTUU婶�6��s�ԩ�������Gt�;����~:���|j������XܞC)pO/z---��>� ���C=      P
N�8��F���r�3fd��UTT���@(][�n�^x!}�� :���؆��^>5bĈ,n�իW�?ݺu��������(m�`���}-F�      ЕR���_�:Μ9\쮻�o~�A��Ci�7o^|��_�q��б�Ѕ��%&�/6l�0q{���J_�i!����?�yTWW      t����\�[��V�y�A>�^���� ������W��_��ѯ_� :���H��Kq�ɓ'��?��O����>� ��w���x����'�      �
�w��>�TEEE���1{�� _RS!p�ҕz�������}�w1�1��E/^��np^mmm���w��A��R�˒%K���.Ə      ЙΝ;���MMM�y)�|��b֬YA���f׮]��6d��}��@��Cؿ̝;78o��Y�ާO���P^ҭ#����㗿��A$      :��O?��:�y)n��c�̙A>i*�<<��s1f̘���hw�d)���~���AD߾}�?�i�ScP~�?�<�L��'?	      �iC�e˂�R�������Ӄ��T@yH7����g���kTWWо���,X۶m"z��?�яb���A����d[�Ϟ=@�X�bEL�6-���      :ҩS��7��M�H����o�����6��o߾x������}	ܡ<x0^x� �����1lذ��ҁL����C��̆�      �#��=��'O�λ����;��/-��֭[�(}/��r�(�_�j �G��$�~���Fccc]eee<���/})(�t���ݻ(/G���s�fCJ      �/^��npޜ9s����!u5)r?|�p ��m(����e�Ў��I��k�֭A��?�ƍ�m�����W_}5�M�f�     �vw���l��͚5+��ޠX��@�;��#G�ĳ�>?�яhw�Ǐ�?���A�]wݕE�P[[@yJ�ǿ��������      �������o���A������'�@yY�lYL�:��Wh'w�O=�T444D�}�k_���/ q��6g������|'      �=���+�u�� bԨQ��c�EEEEP<�B�ICZ��������ߢG���;t���z+֯_E7bĈx���������[�n���@y�7o^L�>=�      p#�9�?�|p����~�}�N1Y���ѣ��?�9����pc�A����?��Qt���GQ]]Ц��2�
�<��?�����       �-m���o~Qt�{��Xt��=(.�;��ŋǔ)S��n��	ܡ����ǏG��W�*���	�T:�	ܡ�mٲ%֬Y�g�      �˖-˾w*�^�z��C�ѳg��ӧO�>}:�򒆶~����/~�7q��:Ⱦ}�bɒ%Qdi�>C��ǐ�<�LL�81z��      p-N�<s�΍���������G��gA�����1����w����CHSXO=�T���D�}��_�������`�p�ԩx���_�     ���ӟ�gϞ�"Ky�5jT@��T�ܹ3��4o޼�>}z6,�k'p��v���_�5v��,p��#p��H���q�q��7      \��7�믿E7gΜ�4iR��4Pޚ����C��g?���k#p�vV__�=�\Ymmm<���>��B�0�~Nҭ@yK����K������      |��������7n\�s�=�J�P�Ғ�5k���ٳ�6whg/��R�8q"��{����OF�=�H�y�۷o�<y2��u��X�n]v�      |��W>|8�lذa�lp�|x�gb	QSS���C;:x�`,^�8����!C�\����!G��l�ĉ�       \ɡC�b�Qd�{���^��2`���֭[455P�N�:�?�|��?��	ܡ=�쳅~��1cFL�4)�Z���m۶�Ǐ�~��      �J���?�������}�{1p���ϒ6����f7����k��]w���rK WG��d˖-�~��(�#F����p�\�����/g����      \(�6l�"�ַ��F�
�"���C�kii���z*����9^����Akkk<��3QT麬'�x"�	�U�6򥡡!�^��?�q      @�����}ERWW�g���
ȏm۶�ڵkc֬Y|15*�����k׮(��~�n���ȧ+V�׿�����[      �ġC���R���#�\-M�˳�>�&M��={���p�������dq�Ѕ�կ_�쥭��>��H��<��s���      'N�����GQu��=�|���ѣG���C�|��G�g�c�=����Z�dI;v,�hРA&�iiJ}�޽��{ｗ=�ƍ      ����s444DQ}�;߉!C�\��STTTdƀ|X�hQ�}��ٟo�	��|��ǅ�.����'�x�d1�"M�!��Νcǎ�~�     @1�ٳ'V�^E5y��8qb��J]N߾}��ɓ�Cccc6�����|6�;܀ę3g�����7��\���k׮x��cʔ)     @1=��3���E4hРx���W��,p�|Y�vm�{�1r�� �L���ԩS�x��(��Çǜ9sڋ��-mq�4iRv�      �����{�ETUUO<�D���Wj*v��@~���������������rw�N/��R���G�t��-{���E��v������;�#      (�����瞋���7�7�|s���T@>m߾=֯_�'O�rw�ǎ�e˖E}�߈�C���t%[�hnn �^|�Ř9sf6(     @1�%H���"���g��Qwȯ46q�Ĩ���b
#���͋���(��n�)n���������Ƒ#Gȧ�G�ƪU����      �/u/��RQϞ=�G�����U[[@><x0֬Y�Ƀ+��5:~�x�\�2�&ȏ>��i1:L�8�C���/�e��     ��k��V��z��߿@{H?K������@����1c�-\�F���/���9s�Đ!C:�+� ��;�]Cy�]w      ������͋";vlL�81���� ���?G��e˖�7�� >%p�k��GŊ+�h�*F�ùR�!mq�={��c     �{�W��ɓQ4}��Gy$�����wȯ�R�q�ѣG� �S�5H$E��2;|UUUt����i�x͚5q�w      �������~���ݻw@{K�;�_i(l�ҥq���p���R�)����ӧ�M7���Ơ8�ϟ��~{6D     @����gϞ����׾�ƍ�����ۂ�{������ҢE�
��=]�u��t��={f?s�O� �:o��f6D     @~�����ŋ�hz��=�P@G�4�/5S���j|���@�W%��-[E��<I�1t�t �C1̛7/�M�     @>���gΜ��y����n�Q����jkkk ����/�׿�u[�!�pU�dTѮ��җ��Ǐ�L)p߹sg ��gϞx���]�     �iy`
܋�+_�JL�4)�#u��=���}�Q ������k�o}+�������
w}VUUU|��ߵU�N�J-(�����     rbɒ%���ޭ[�x��:Cj*�,ȶ���(2�;|�U�Vŉ'�HfΜ)4�K���bI�ӭ#G�      �Wccc�&w�}w���t��Tl۶-�|;y�d�\�2�瞀"���hmm-��Y555�t�;ϢE������     ��|��,�+���y���0�cΜ9QYYPTw��6m����G��{�ѳgπ�п��z�s��P�֭�����_80      (?---�[�<��ѭ���ci Ǒ#G�7ވ�3g��,�E;�6,�L��U***����@��_x�����c�      ����_�ÇG�����m��Й�P,/��r̘1#멠���<�mp/���ߵ&t�t �C������=z      �e�Q$UUUq�}�t��}�fߩ644�{�쉍7�����H��!moomm����W��F�
�j&��xΞ=k֬�9s�      �#�w�w�"����cРA�-mq����}��Pi���������n���Q���{�(w(�ŋ��w��j-     �2��IMMM�u�]]E�Ųe˖صkW|�K_
(�;\��U�
u�ϤI�bذa�@�Ŵ������E      (}�M�6E��s�=ѳgπ�����Y�ti���?(�;\���ˣ(�u����7JE�6������� ���W_�     ��E�EkkkE
��N�Е�P<k׮��<���P$w���͛u��̙3����"]0 �;@����[q�ĉ��       J�ٳgc͚5Q$�������*�+	ܡx���������w�D��HE�B��o�=�Ԥ-�w(����X�jU<���     @�Z�lY444DQ�9�MĔ��STVVFKKK ő��x ����B�8y�d����Q3f̈�}������|@���kq���g��     �����H�+**���P
�2�~��e7c�q�ԩX�n]̞=;�(�p�+Vd�c���vJY�8�)�ްiӦ?~|      Pz6l�G����4iR�1"�T��_���
(-�S$w�?����r��(�iӦe�P��a(�4p&p     (ME�ޞ��{��$5[�n�X�m��w�[n�%���ҋߡC�����;�(Uw(�w�y'�^�o߾     @�h���(,�i*���-[?���@���H�ۧL�� FI����޽{�ٳg(����x���m�      (1i{{KKK�偔���� �i�����ODϞ=�N�����!�|��(���*0�B�8���(��˗�     JHZRdy t=ܡ�R�v�ژ3gN@�	�����Q__E�`(uw(��{���ݻ�[n	      �������ɓQ�R����mo.J�\,-�Sw�_�V��"p ���8��'�|2      �zE��>y�d�)i�����0�xv��{�쉛o�9 ������c�֭Q'N����;�����������      �Ή'bӦMQiy�]w�P�RS!p��J}SOy&p��֮]���Q�g�(w�ԩS�y��7n\      �uV�^---Q�R�w��R����G�n`��O7���"=zt:4�\����KXSSS ŕ>��      ]+�tE�n���r`i ۙ3g��wߍ)S����Bۿ�ٳ'�`֬Y�$�� M<x0��z��7�?�aTWW      �o۶mq���(����flʁ�X�r���\�Shk֬�"H��o��r�dw(����l�x�ԩ     @�[�zu��픓A�e?�---ӆ�ԩSѷo߀<�Sh���zA�ޞ^j�ܘ8��y-p     �|���ٍ�E0v�X�QS6�u�-�<v�X Ŕ\֭[��sO@	�)�]�vő#G"�w��*ʖ�߀$M744D�=     �γq��8}�t���PN�@���--��Ww
뭷ފ"�<yr���3����s��e�<��     �s�]�6�ছn�[n�%����b˖-׶m���ѣ���Kw
��{EEE̘1#�\��X�9nmm���՗w     �Γn�}�w��㎀r#hRS���?��y#p����������(Wݻw�~���G}@����������     @�{���=��ƍ(7ii �����SHil̚5+�ܥ��������{/&N�      t�7�x#�`�̙QYYPn�@�gϞؿ>< O�R�2λt�J�����QUUP�ҁl۶m��[o	�     :A���K�O�<9����D�^���?��RO!p'o����ǳ���kii�g�y&���ƦM�(7&��6��n���FEEE      �q�y�hll������޽{���T�޽;�b{��7㡇
��;��~��,�+�ӧO����cŊ1jԨ,t7n��(w�ͩS�bǎ1z��      ��M�E0cƌ�rV[[+p��>���;����Q���oߞ=}���I�&e�����2�;p��9.p     �8is��"�7�tS@9�T m�pڷ��퀼�S(�Ν�-[�Dѥ���S.�@FϞ=���> R��裏      c�ƍ���y�������M>E��m�|�M�;���By���ȝ�.��>hР�:ujL�2%jjjJI:��ٳ' ҵZG�ͮ�     ������Q)ܴiS�����ٳc�������@��;wƉ'b��y p�P��W��رc�hѢX�dI�;6�Ꞷ�WTTt5�;p��5dΜ9     @�J���w1E�n_�n]��F"������
(i�e�ymnn���g��⮻�
��;��6����o:��'Eœ'O�6����;���8.�6i�     �ߎ;��ɓQ4)
ܾ}{����7&M�ӧO�������s�n�H������8t�P9r$�z�?���}�ҥ1f̘lRy�����Up��6o�---QYY      ���ݩS�b���bŊO���7�wS����R�$ipcccTWW�;�;����r}���>��B�4�<eʔ�޽{@gH�1�6gϞ��;w�     hg��Npޅ[�S�N�Z�����R����$���!�l�uuu�N�Na��$n��Çc޼y�x��?~|̘1#�Б�]���� I�\�     ���Ǐ�޽{��;v,-ZK�.�1c�d[�}WE�����6�6�;y p�ZZZ��$�O��Z�n]��1";�M�8��&t�����ȑ#�����      �ǆ���|����ظqc���ٓ'O�z�^�zt����&��7P���Ν;��ٳA�طo_�,\�0���5kV2$�=���h��������={      7nӦM��K�_���˖-����ǌ3bذa�m����&}>����N�N!l޼9�x)4�p�{
��!.m߆��Pssslݺ5��     �ƴ��h+�SCC�E�D��>q�Ĩ�����޽{[�	|"�͙3'��	�)�>� �\i��ܹs���mWr80�z	܁K��w�;     ������̙3��I�DzR+QWW�-2dH@GKME�s����{wʞ���KS�۶m���ӧc���bŊ5jT��7.*++�����6     ���6��~���?��~뭷f��رc���*�#܁����Y7�ѣ�	�ɽ��t����ؾ}{����7&M�3f̈���\�����v�ܙ]�أG�      ���M�t�ԭ��O�>1y��>}z0 �=���@��g�fM��ѣʕ���۲eKPZN�:�mu_�re�9�Vw�J
X�pD��H���cǎٶ      �Ϲs�eut�ӧOg�Ċ+bԨQZ	�U��p���]�N9��{|�AP��5(m[�S�N�)S�DMMM������P���     \���}SSS�9Z[[��;�;p�����
(Wwr-
�m���cǎŢE�bɒ%Y��&���rEEE@�t Kۚ�lݺ5      �~v��e���ѭ[7�*�'� UsssTUU�#�;�v���8s�LP>҇�ƍ�'�̓'OΦ�{��`���Ν;�A\�     p}҆W�֕Z�����+�j��KS�Z)����!>���lp
ʑ��\KSH��#G�d��K�.�1c�d��ѣG�%p.U__��n�)      �6i۳[�K˅�D]]]̞=;��ERS!p.����+�;����@�6�<bĈ,t�0aBt��=(�;p%i�M�     p�RW������J�_�>{�Z��'Fuuu�������>�������ʑ��\��Ͼ}��g��1~���1cF6,(�~��e��Ν�6�����      ��֭[����J,\�0��>k֬2dH��,.�>�[[[���"���ɭ4a�w�� �bݺu�cR�8��V�8޿ �1�     p}�m������OZ�[o�5�ǎUUUw�R�q�Y��ʍ���ڽ{wv]�gR�XҁL�\(���~�׳g�      ���ܹ3(O~�a����'&O�ӧO��%p�$-�S���֮]��b�pR9}(��}���&�sƁ�T�NkϞ=�|%      �:��S�N����ӱ|��X�bE�5*�M��ƍ���ʠX�B�4�~& ڤ���;�(7wr+mp���F��s�f[�Ӥr:�80(w�J���     ��m߾=ȏ�*�w��~���ԩScƌQSSGmm�����{ʕ���J�0�I���Wb�     �ڤ����ɓ'c�ҥ�lٲ;vl�J�f���"ȷ�T�ڵ+ ڤE�����-PN��RSSS�߿?�ͅ��}���I�&e������K�6N
---��`     ��ٹsg�o��ͱq���I���ɓ�ؽW�^A>Y\*us�3?<A9��K)nO�;\ɩS����+W���#G��ٳ��n3�\&�u��cǎ@�����w      �/��{��	��ȑ#�hѢl�{]]]�J><��;p%�f�;�FD.�޽;����m[�S�N�)S�DMMMP�ҁL�\����[n�%      �|�{���Ơx��j�ׯϞ#Fd�'L�ݻw�_mmm \JOI9��K{���)�n�T3fLv�5j���%*�[�l	��۷O�     p>��À��Zz.\�mu�5kV2$(_�n�N� m|�S���R�4��^�7nܘ=)��<yr����+(�����?     �ձɕ���Ǻu�'muO����㣪�*(/i��A��СC�&�����=z�(wr)M�:r��e[�G�t=�;p%>�     ����ϒ�s�;wn��=-�>}z0 (���jmm�={�ė���r!p'wҤщ'�˅[�Ӥr
�'L�ݻw�����     �X���|�ӧO����cŊ1jԨ��7n\TVV�MS\I���SN��N�$M�1���+=,Ȯ�1cF6,�\�{�Ξ�g�@�ÇGcccTWW      W�n3������پ}{����/�N���555Ai����K��PN���t�tS��u벧m��ĉE��h����k׮ h�~�v�����[     �+KK��z�<y2�.]˖-��c�f�D��^QQ�܁+�URn��N
۠3�mu_�pa���ŬY�bȐ!A�J2�;p)�;     ���q����c�ƍٓ���<yr����+�z鿓4t���1�F���;�
�
�
�����zk���媪����R��Ç      �M�N{:r�H,Z�(��>f̘�={��T]�G�ѧO�8u�T �9{�l|��Gѿ��r p'w�m��?�0{���S�L�&��ܸt�َ;b�޽�?\�{      �������>��>bĈ���0aBt��=�|i����TzаQ.��J�ZG�F)I���^{-�/_��v[v�K������;v,�y�x�������y��     ��RW�{W:ھ}��g�QWW�f͊!C��'��J7�;6��ɕt�FCCC@�iii�͛7gπb�ԩٓ���r�*�?�U�VŮ]��j	�     >�ѣGut����X�n]����)t?~|TUU���6 .�ʉ��\���rp�ĉX�xq����D\��>j�([��|ؾiӦX�dI9r$ ��ɓ'�_����3      �����B�<w��l���ɓc���ق@:F��p)K)'wrE�N9inn��7fO��M�{:����;�(f_z�ػwo ܈4 s��7      �U��N�>˗/��+W�m�ݖ��_��W,l'�q��yǎp)���;�r�ر�r���[�`A�ٽ��.��o���(�������իWGKKK ܨ�w��     �r�6JE�6oޜ=�:�)S�DMMMpm�����~l۶-8���p%��lll����R'p'W{�_�>{��M*O�81z��y��,?����0@{9~�x      p�C�����ޢE�bɒ%1nܸ��9rd��Μ9o��F֗襀��`R�5|���R'p'Wm����㥗^��_~9ƌ�f���V�49���OG}}} �'��     �2�)e��ͱaÆ�<xp�O�4)z�����G�k�����i�"��J�wʁ��\��G�@�q���馛���������u��e�~�r��	�     .׶��A
0�͛���J�H�VbĈQT�t��x��ׅ��1�F���+w�n�޽�3��� 7s��:th����z+^|���' ��      �������ƀrr�ܹx��7�'/K��{���_�ԩSp���;�q��٨��(�4�����'M(O�6-&N�X���?����v�C��     p9ߡP���Z�����~����^,�\�ɍ4iE�o߾�I��)S�d���A��Լ����v�S�w��wMEEE      p����h[
����92��>v�ب����H���ٴ�;���;�!p���-+V���+WƨQ��нTp{��^xA�t������Ě��      �<[ɛ� �ر#{�����R�D9���������<ڛ�ʅ���8u�T �p۷oϞt��<yr6��U�3g�ğ���,8�,'O��     \@�F��>}:�-[˗/�d)�q㢲�2�I���z�8w�\ t��Y��c�w�P���F
ـ��\:����]q�K��s�=��'��ҁl���     �yǎȻ��E���H��ӂ�R�u��ls{SSS t�4�6t�ЀR&p'7lp���U�%K�Ķm����     �؉'�$�̿��+�t��;vl�J��Qj����ӟ��@��S�䆐�N�.���v[̚5�Cp��6�t�      �ST��ͱq��쩭��N�:5z���������SOŹs��3|��G�N�Nn��צ��%6oޜ=�}�K��͛����     �������ѣ�hѢl���1c���G��?��x����:���r p'7Μ9��i�����cǎ�U�      |��ٳ����yMMM�lu1bD�IL�0!�w�ީ�>R��k׮ �L'O�(uwr#ƀs�n�С1}���8qb�����5���c�Е�      |ʦV�l���˞�:L�4)k%���w7o��V�
��潀r p'7�lо</��R����QWW�gώ�Ç�?o͚56']��?      γ��XZ藚���muOK������VCCC������ ��{�@�Nnܡc����ׯϞ/��+]i�v�� �j�      >eS+\����K�,�ɓ'g������_�ҥ�\]��?��;������ �`��?~|̜93������7ް�(	w     �O�>}:�k���,_�<V�X�F��B�q��Eee�u�k>|��@�K	�)wrA��+]��nݺ�i��^WW�W��R��      �S���imm��۷gO߾}cҤI1cƌ�߿�5�k��/���� �*�
ʁ��\����k�mu�?�������      ����O�|����Z�*ƎӧO��#GFEE��s�n�;v�����������m����¹s��Z�v��455e[��H      ygS+����}�ƍ�S[[S�L��S�F�޽?�bŊ �j��H�o555�J�N.����X��޽{      ��б�=�-��K�Ƙ1cbڴi1z���w���g{;P2����R&p'� ������      �̙3t�t�t�V��Ç����c	���+W��R�vJ���\� ��~      p�������/��B,\�0���bӦMP*�P��䂀 �Tccc      ���@ר���u��@)�n@���w �R�      ��	 p!��:�;����  ��     �< p!��:�;����  jmm      Dl �żP��䂀 �Tsss      ��[ �bwJ���\�� ���     ����&ߛ  �S��䂃 p)�      6 �rnw��	�� p)�      �3 .���P���� p)�      �3 .���P���BEEE  \��     �� ���:�;�PYY  �~      `C+ p9p�:�;� ` .��      ��V �rwJ���\� ����
     ��� ��~@���w �R       ��Z[[J���\� ���     @S \���N�N.� �K9�     �� ����R'p'�u� \�{��     Pt6 �R�(u�`rA� \��     �� ���J���\� ����     ��� ��~@���w �R�      l �媪�J���\� ��~      ѭ�< ����R��\� J�H�      "��� �B�KJ���\�ѣG  ��ٳg      p~1P�����  ���R'p'z��  m�      |*Elw ����R'p'��4q���  w     �O����ٳ ��)uwr���"z��gΜ	  �;     ��Dl �����J����H!�� H��      �	��y7��	���Z�6�      >e9 p!]�N�Nn8� m�      |J� \HWA���}�� ��_�~     �y"6 �B��(uwrC� �1�     �) p!��:�;�!d �|     ��� hӭ[��޽{@)��B6 ���7     �O���+  ���;�!d �|     �TMMM  $nv���! ЦO�>     �y�
 �M���J�����. ��I����      ༾}� @⽀r p'7R�^YY--- נA�     �O�� ��^@9��)nO����� (.�;     ��Ҧ֊��hmm ��lp��ɕ�
����      ����޽{Ǚ3g (6�)wr%m۷o ����      K1�� ���r p'Wm ��     ��0 ��� @��*(wr�_� ��     ��� ����y��u�����0�0�30ð�"��b�7�D��W�TJ��m;��{�U7�][��ʹ�̫�l�i'��Ina*����2��,2���t��PYf�.��9�3�R�����|>���xO@>�SP (n���     �_�իW  ŭ[�nQSS���A ����l{M      ��i� @z?PRR����������  �O�{      ��� ���B�NAi�ںq��  ���\      vM� x?@��Sp���#p�"%p     �5[ ��w
N
����? P|�      �VYY555�y��  ����|!p��� (NMMM     ����B� �K_I��Sp��� @q�>      �ͥ���V�
 �8	��w
�� �SUUU���      ��w �8UTTDMMM@>�Spz�oݺ5 ��a�     �[3� �WZ�VRR����ܷo�xꩧ (���      ޜ� ���\�'w
R��*p��b�;     �[K������  ����|"p� ��
 �ǅ     �[�������ظqc  �EWA>�S���� (.��      o/�@�18�|"p� 4( ��&����      o-Mo}�� (�������/�����,tkii	 ��80      x{)p �KCCC�����;+Mq�@q�     ��; ������;+�n<�@  �O�     �{R�VRR��� �;�F�N��@�H;�      ��z����/ P����;k��� �����ݻw      �{R�&p��ap �F�N��իW���EKKK  �k�С�6�      ���w�} ���J��;w
Z
�V�X @�J�{      v�)� P<�y��@����&p��'p     �3w (�7w
�� 
[Za�|     �gjjj���.ZZZ (lw����6dȐ(--��;w Px���UUU     ��IM��~��  
����#�;�{��1`��X�fM  ��E     ��I�Y� P��������|#p���9R� *��     �sÆ ���m%%%�F�N�K��w� @�5jT      ������s��  
S
�!	�)x)pO+�Z[[ (������      칊���߿�]�6 ��d�����WSS}���u�� P8Lo     �7i��� 
S<dȐ�|$p�(�)�w (,��     ��1bD�� ��������H�NQH^�_ P8�      ��� (\���|%p�(�3&�n���5 ��WWW��4     `����;;^|��  
��l�3�;Ea�������X�fM  �o�ر     ��K�� 
���|&p�h�)�w (w     �����˗ P8���uuu�J�N�H!��� @~+))�ѣG      ��tW (<���;�;EcĈQ^^۷o  577GMMM      ���	�--- ����? �	�))nO��ʕ+ �_iW      �Ϙ1c�W��U  ����$F��������� ϥ�9      �G� �c��ѳgπ|&p��p�q�7 ��z��Ç      �O�A7M{mmm  ���k�������hjj��> ��������      ��&���v��  ���B p��L�81~� �&L�      ��4�]� ����<F������	� ����f�     h)p���� �_#F���ݻ�;�;E'�N����-[� �?����     @�5jT���#^}��  �S �@�N�i����_�: ��1q��      �c���Ř1c���  ?	�)w���,p�<���      t��	� ?���/���P��q��EEEElݺ5 ��7hРhhh      :N
�KJJ���5 ��bz;�D�NQ�޽{�[u ���v     ��WSSC��'�x" ��"p���)Z)��@~8蠃     ��7q�D�; 䙪��>|x@��S��Yyyyl߾= ��5`���۷o      �����[n�% ��q�DYYY@��S�***bܸq���. �ܕn�     �9����_�~�nݺ  򃶂B#p��r�!w �qS�L	      :O��~�� ��*++c̘1�D�NQK�r���#^}��  r�СC�O�>     @��@��0aB����;E-����}��� 䞴�
      ����9B�~��  r[Z��F�Nћ2e�� rPIIIL�4)      �|tP�v�m ��ݻǸq�
����7f̘����M�6 �;F�uuu     @�K;�
� �p�QQQPh�������?�i  �c�ԩ     @�8p`���?�}��  rӔ)S
����a�&p��V|��     @�I���� �{���b�ر�H��k��1hРx�� �z�'O��     @KSao���hmm  ����[70��o6���ӧ� G��U      �Z1t��x�' �-i�(Tw�?i����Ŏ; �:MMM1lذ      �륞B� ����>F�P������������ t���JIII      ����3m�4mM�o0c��; t�����"     �ܐN�81��  r���B'p�7=zt455���? @�;�����.      �i^�; 䆑#GF߾}
��� m�q���M7� @�{�;�      �q��E}}}lܸ1 ����A����8����[o��۷ �yc���      rKiiiL�2%n��  �NEEE|���N����:&M�˗/ ����i7      rOx��Gkkk  ]c���QYYP��)��@�)//��     @kjj�Q�F����  ��GP�Æ�!C���ի �xiK˴�
      �+Euw ����Y��@�o��|g|��_ ���.      ������hii	 �s͜93�X��ML�<9n��fe ��ƌ��2      ���������G?�Q  ����29䐀b!p�7�.���Z��zk  ��v     ���Z���Ǳs��  :ǴiӲ�����B�(�����ؾ}{  �O�>1a       ?���g�w���  :Gj����-���Ĕ)S⮻�
 �����%%%     @�H�x� �9ƌ(&wx�gώ��;Z[[ h?���1}��       ��=:���c�ڵ t�#�<2����m455Ł+V� �������       ��)��^{m  �O�>1~���b#p�����w hG)l�9sf      ���N���rKlڴ) ��������;�!C�ĨQ���G `�͘1#���     ��ԭ[�����  �_UUUz��H��)Mq���+++�V     ��Ҏ���~{l߾= ����UTT#�;즱c����c͚5 콴]e�^�     ��V[[�M���/~ @�I;�H1��n*))��s��W���  �Niii�+
      �a���q�w�Ν; hӧO��={+�;�<0���c�ڵ �iӦESSS      P����{�7 �}��}���L�{ Mq�7o�)� �Lo     (L�z׻ⷿ�m��� �o�±>}�3�;�!S�`�L�2��v     ��:�ѣG�ʕ+ �7�sL@���JS��ΝW\qE  �'Mo�3gN      P��=�X�; �������������A�5k� ���M�fz;     @>|x�5*}��  ����'w�i������K_�R  o�[�n��'      �4��s��\  {nܸqق1@�{-mb�1 ��#�8"     �:
- ����/���K.�$ �]����w��]     @qH;�
�`ό;6F����a��@&L�>�`  ��#�����      �8�=:F��=�X  �g޼y����Q����CEkkk  Q]]�sL      P\�?����K x{'N̆�!p�}����zh�}�� �EZ]ܣG�      ���Ho	��� ��JJJ���~w M���㎋�����u��  "�#�      �S����CEkkk  �v�!�����kwhuuuq��G�~��  "N<�����[M     �b5`���<yr��7�	 ��ű���SA;�={v�u�]�q�� �b6jԨ8��     ��6��X�bE�ر# ��v�a�E�>}�{wh'ݻw�VS]{� Ū��$.\      ����~x���? �/***b�ܹ���ѡ��]�=��� �(�      �̛7/��x��W ��c�9&����5�;�����X�hQ\r�%��� PL*++�m&     �MMMM��]o�9 ������>:�7'p�v6lذ�:uj,_�< �����={      �ёG���/�^ (vix`EEE oN�`��q����^��ѯ_��9sf      ���֭[w�qq�UW ��ƴi�xkw� ���1gΜ�馛 ��I'�eee      �2y����OO>�d @�:�����$��&p���׺��cݺu �,݌;vl      ��I1ߢE��3��L��� �I�&�������CISl/^����\�P�*++���      �vӧO���+ �����ǂ�=w�@#G�ta@A;��㣮�.      `w��K+V��-[� �9s�D�޽�=w�`i��<�7o ($C��#�8"      `w���ļy����n @1hhh���>:��'p�V]].����: �P���Ʃ���}     �=1k֬���c�ڵ ���O���� v��:�ԩS�W��U<��# �ਣ���      �4DiѢEq饗Fkkk @�?~|L�81�=#p�NPRR��vZ�˿�Klݺ5  ����Ҷ�      ��F��vX�y� ��{��ق.`�	ܡ����;�ϟ7�pC @�J���8㌨��      �'�pB����y�� �Bs�q�eC�='p�N4k֬����� �G3gΌ�#G      ����X�pa\}�� ����9���#p�N���.Y�$>��O���� �I�n$      �^�M�˗/��+W ��	.^�8����;w�dMMM��w�;n�� �|�v�UYY      О���d��m� �����aÆ�����:�x���� �3f̈q��      ��>}��q�7�xc @>�ݻw̟??�}#p�.PZZg�}v���klٲ%  �544Ă      :ʑG+V���<  ���Ē%K���"�}#p�.R__��̮�� �\ն(���2      ���(��N�O~�}�� �|3cƌ3fL �N�]�����S��=�� ���̙Æ      �hMMM1o޼����� �|RWW�| �C�]lѢE�jժذaC @.4hP�     @g9�cbŊ�z�� �|�v!Y�dITUU�>���z��g�uV\z饱s�� �\PQQK�.����      ��RZZ�=������k�� ��f̘�Ǐ���!><�����   �r�)��      ��c��o}+  �544Ăh_w�s�΍������O t�I�&����      �J����#�Ľ�� ��Ү#g�}vTVVо�#�Nv���'m�@�I+��,Y      ��/^�V���7 �9s�İa�hw�!)*<���k�	 �lm��z��      �ժ�����O�/|���� �+��@��C��>}z���=�� Й�?�x+�     �)cƌ���:*~� 䂊��l�`YYY C�9hɒ%�nݺx�� :�ĉ�裏      �5���φ�Y�& ����=�� :��rPyyy��}�O}�S��+� t�޽{�g�%%%      ��[�n٤�O�ӱm۶ ��2y��6mZ K�9*ņ�sN|�_��;w t��EU���      ��_�~�`������ �cɒ%t<�;�1c�Ĝ9s�?�A @G8�SbРA      ���xG<����� t���HX[YY@��C��7o^<��S��� ���;,?��      �|PRRg�yf|�ӟ�^x! ���x�1x�� :��r\�8;묳�3��L�_�> �=6,���      䓪��x������gc۶m m���1s�� :����/ζn� �/jkk��s�Ͷ�     �|�����zj|��_ �HMMM�dɒ :��	�Ā��UW] ����ʲ����>       _M�:5�x���� �***������t.�;�C9$�8��; �ƢE�b�ȑ      ���O�5k�ĪU� ���ŋ���t>�;䙅Ƴ�>�<�H ���5kV̘1#      �t��-����O}*ZZZ ��QG��t�;䙲��8��ⳟ�l���7n\�t�I      ����6�=�������رcG ��=zt,X� ��#p�<TYY\pA�ۿ�[l޼9 ����/�9�(--      (4Ç�N8!���� �޽{�ҥK5���m�.��2+�xS��_�(�G�      ���#��5k�į~�� ��Q^^�}�{���&��%p�<6bĈX�xq\s�5 +]x-[�,      
ݢE���}�ڵ {���$N?��<xp ]O�yn�����K/����� �6��묳Ί�C�      ����x������g���% `w͛7/9� r��
@:�n޼9~�� $'�tR|��      Ť��.�?�����Kc۶m ogҤI1w�� r��
��'�7n���? (n�gώw��      �h���q�gƕW^��� ofȐ!q�gDIII �C����4�.]�]vY<��@qJ�e��      �,�v|��ƭ�� �+�{��.� �w�@n�CI'ڴ�ֿ������? �1c�XU      �gΜ9�~��X�|y �UUUŲeˢ��6��#p�SSS����K/�6 �aذaq�y�E�n��     @�C�v�i�y��x�� ��V���������PP����㢋.�"���� ��80����GEEE       QVV�{n|�s����~: (nm��F�@��C�jll�}�CY�iӦ �0555�>��l�,      ��UVVf��.��X�~} P�.\S�N �	ܡ�����/�V!oٲ% (,}��/�8jkk      xs555ٮ�)r߼ys P|fΜGuT �O����9�@���?[�n 
C}}}\t�Eѳg�       �^ �lٲ�����^ �G��~�)���P��~\~��}��  ���)n�ݻw       �oȐ!�| ���/P$<��8�3���$�� p�"1z��,r��;v� �SUUU\x�ѷo�       ���������j( 
ۘ1c�sΉ��� ����رcc�ҥq�W�Ν;��RYY�Mn8p`       {�-x��+4 �mAS�nRY�7��B�9蠃���O�k���@Iq{�*q���      �<0�8㌸�ꫣ��5 (C��:���� ���дiӲUi_������_ r[UUU����aÆ      �~�N����^{���@477g�E&�'�;�ɓ'g'�~���}��  7����E]�]|      �o�����k��7� �>}�ą^����/�;����g۰|��_�.� �-={�������      �q���wƖ-[����~ ��z��u����7�;�Q�F�?��������J �z�>766   �-�رc��}�{���  @~�7o^l߾=~�� ����..��⬷ ���!C�d+׾��/��/� t��}�f�����  @�Ν;�)z)"O1y�ұu���{���j�1}���g?���?���f?�>�}�~����+�L:v���RRR��<�����]}��������O����ʲ�����\^^���+**������ا寧m�Zڞ9}���
   �����]��v�m@~HQ{�,(w 3hР�������?---@�8p`\x�QSS   �b۶m�y��?��)VOQz:R�����������):o;
͞��)�o���t�ħ�-�O1|����6��G�QYY�}La|:z�����  ���p�	����o�9 �m)j��?(n���3�g������q�e�ņ�Εv���>��,  �Ui�?��Y���+�d��H�-To��S��>���s���.$H�wW����I��c[���t��b����/�ӑ�  ��fϞ�����|ǵ-@�J�[��^WW@a�%�d��⋳�}���@�5jT\p���  �Ζ"��7f��7mڔ}�"�4a�m��`�]i�}H��ۤߛ��65>M�O�H���t�§k����,�����~  �+̜93[�{�u׹�1��/�0���;�wz��Mr����㩧�
 :�Ag�}v�0  �=�����HS�����i�)H��UڦƧ�����V�b�tݜ�����)�Oӹ��� ��2cƌ��ꫯ���F�˖-�& �I��Rz8�&����g���@ǘ5kV�|����  `w�M]O�_z�l�z�����q�6�7���w<���J���"�4>�'555ّ�u655Euuu   �C9$�ָ��+�]� �:�F��.���(pw�M������}q�-��m�� ���ϝ;7�=��   �[)�}��c���Y̛&��p�m�q���ߋt��'iǂ�������S߽{���g������eccc���  ���8qb�w�y�|E��E&L��}�{�!@a�o)m�{�	'dx����lR ��[�nq��ǔ)S  (^)T߰aC��	�i{[��A9�����?�n�����#�<��_�L������uuuY ��ܜ��  @q7n\\x�q��g�� t�ɓ'�Yg��ݿ
���-3f�Ȧ]u�U�m۶ `龜�iw��e  P�^~��l
{���D��y
kS��	���o����Y����{���o߾��  ��0r�ȸ袋�K_�R�� ����ŋg�Z�� pv���G���i� {&톱lٲ��7  P8R��nݺ,do�طnݚM��C�x��==\M�{eee���D}}}455e���  Px���ǲ���� :��ٳ��㏏��� ����#i+ޏ~���E�ڵk��3|��8���  @~j�ƞ\��5}�B���-�Ȑ��#-tI�N|���{m����o�l�{�>}b���Y  �4�*	��W��=�X о�@�E��G@��{,=����?W^ye<����[�>}z�UV�n�z @>x�����"���]
ٷmۖ� {ꍓ�7l��?�x�}���C�4ݽ��*jkk��}����W   ?TWW�E]���7�7��M �>***b�ҥ1q�� ���
�+i�������w◿�e ��҃�M�1�  @nI�z�ľnݺ,dO�_}��,d��u(E��H�C�W�ξ��'���)|�ٳg444D������>  �ܓ�\�}���{��o�= �7i�\C�	�x	܁��.�N=��l;���ر# ��4�!�&;vl   ]+E�)f_�vm����iӦؾ}{���@�I�{Zp�����O<��雷��!occc6�}РAv� �PRR,��}��u�]�����K���-[�{�����	�3fdo.��կf��]�q�v�hjj
  �s������3�ĳ�>�MD~�W���bv��;6lȎ�+Wf_K�{Zh��E�E�555  t��;,z���i�& v_ x��F�=@����Ç�'>��"��'��b5q��l����   :N�p�~��x����---ٴ��u�b�v������W��_���QZZ�ݛ�������)~O_  :֘1c������/����Ҁ�E�EYYY $w�ݤ�%_|q|��ߎ��+ �Iz@<��8�c�- ���&�=��ӱnݺظqc6�=M1`��b�-[�dG��"I�+***���6��{���!z ����k�E�k׮ v-ݗ8餓b֬Y�Fw�]����i���F��믿>�n� �.m�����i  ��IQ�3�<�=�}�bӦM�}��hmm �^zM�ґv�X�re��{�)zoll�"��  �������h|�[ߊ�˗ ���:�9���Kw�CL�6-W\qE6]�P�92���ٳg   {��_�5k����?---ٴa1;@�H��iG�6dG�������l�Φ��>|x��  �siA�g�����[n�%[�@Dsss�w�y��� �"p:L�~�������7��{��B�&��-�.\eee  �������g��B�W^yŃ]��^���u:����+�{��_6�2�9C���ݻ  ���s�ٳgg1�UW]���(f�'O��N;-***��܁�&����&L�뮻.����Բ�O?={m  v-��<�L�]�6�ξiӦx���Mg�C�����cv�^�:����֭[���fS��i�;  �k�ƍˆ~�+_�u��@�I��ϟ�sL���܁N1mڴ<xp|�k_�n�ѣGǙg��m�  �EKKK�Z�*���H��
ێ;⥗^ʎ�+Wf�{��My4hP6̔w  �i��'>�����w�uW �4H�Ί�c������_�~�},n����; ����s�̉y��YI  ���_�'�x"�8����۷{�P��[�lɎ��i���Q^^�MyO������a6  ��>���N�Q�Fŷ����
@!9rd,]�� A`�܁N�.�N>��1bDv��v ����8��c�С  ��瞋'�|2��&����� o%�:iAT:~��(++�"�4�r����=  (VӦM�����W\6l�B��̚5+.\�� �w�KL�4)[�w�5��C= �*�XZ�hQTVV  ��;w��ի㩧��^x!^~��l2/ �tٱcGlܸ1;y��Awuuu���7���=i=  (������o|#x�� (UUUq�g� {C�t��5�e���;�o�1�n� �"M[�d��-  ��k�����O?�t6e7�&h���sMZD���gG
�{���{�����l�{�ne P�Ң���??k'n��l'$�|6t��X�ti444��rW�R�Ō3bĈq��Wg��ڸq����O��={  �m۶ţ�>�]����K�� ��R�Y�c͚5�|��lW����6lX6�҄w  
Q[;�y~�k_�g�}6 �Mz-�5kV,\�0���`_܁�Я_���G>?�я��?�q�U-@gK[d�x�1}��  �B�s��X�zu�Z�*^x�x��W r]
��9+�0����<M��۷o�92���  
I������x�|��q�w@�������>;�^hw g��{�{lL�4)�����;@g?~|�z��E  ��{.{�X�n]����Y$ �,���9���ώ4�}����>}�Ę1c�w��  ����<N>��l����_���J ��z-^�8[��^�@�I+��4����gq�-��&�Pij�	'��m�  ����%�׮]��9Mm�B��u�6mʎ��gϞ1`��;vlv�  ���ɓcԨQq��ƃ> ����2.\�� :���I�AđG�=���7��m����M�SN9%jjj  ��k����|O=�T��⋱}�� �b����7f�C=�M�L��<8�"�{��  ����6.������;��o��[�@.H�L�y���� A��~��Ň?���{�������v����-����  �;vd�W�^��h�[K��֯_���{o6ѽO�>1bĈl�;  䃒��l:rZ�y��Wg�� �JZL>��lpiz}�(w �7CӦM˦��t�M�|�� �iw��3gf[  ����%��Ӕ�M�6Ekkk  {.�C� �'�|2;��ʲi�)tOCҶ�  �������G�g?�Y|�{�3� �tÆ��N;-X
���@�H��6ӧO�뮻.��� �]��SO=5ے  r�Ν;�)\�V�ʮ{�m�&j�����ƍ�㡇���7���  �4�+MM�8qb\{��裏@GKSۏ=��8�裳�!�� p���������w�qG���?�*xK���1w�ܘ5k�-  r�k��+W�����	����q:�#�C����&Ӎ92�w�  �KҢ�}�Cq�wƍ7ި� :̈#���MMMЙ�@^J+gϞS�L�[n�%�/_ o�Dv�a1���o��  r�s�=�E��֭�W_}5 �ܑvTy�����{�=zD���c�رѫW�  �\PRR3f̈ѣG���_������TUUł��"�� t6�;����3�<3=�и���g��Q���;}������Ir��@¾( ⾡�(�-ڷ��u{z��{k��<�5U��>������wf����]^���Kk7����l�����dO���"\�n[� Y^/�S�sN�]b��������]���/bٲe  S���H�2��ѣq� `�K;���Ç�TTT��ʕ+�;�c   7]js������O���������C<��C���Q__ 7��;0#������x�w�W^�7��g������<_l �ͦ� f����hooϓ������˗�]wݕ��  �f���{c͚5���/��o��k|)s�w�w��fpf�Ԝ�e˖x����^�m۶��̗n��_�U���?����  ����ɓq���8w�\ 0s��Pooo�۷/O�X�%K��}�ݗw �-�7M;]�_�>������� �&�,�y�x��d.�)C��q�[jp~����׿�u�޽��d���Л6m������5  7���D?~<:�C�Z��522��Z[[s!KKKKn�[�ti  ���z���?���Ď;b�֭��� �w���?��X�hQ L%����`���������/⥗^�#G�03���Ń>���.  ��R�=]k<x0:::,� �&������ӧ�{SSS�~��  7B���aÆ��{����w�ɟk$)W������{�7 �"w`ƻ��������y���q�ĉ ���z����+W�  �QR#�}������^�v ���^��������X�vm��:�P  �S]]]����a�_��q��� f����x��b˖-yA6�T�;0k�P���_�+v��������`����[�g?�Y�[�.  �FH[7��q������ �*5fvvv�����>����X�jU�y�Q,  ��T �?����O>�$����3!0{�]}�������FCCC Lu����N�z衸�����W_}�ELq��rK������y  p�uww��Z[[��ŋ p��a��0�q�ݻ77k.[�,o_[[  p=��ʹ���wߍ������ f�T
���ݿ�ל Ӆ�;0+�����?7n�?�0^y���0Ť��-փ>��  ��r�,;u�T��� �����i�����s�=5�����  L����x���G�!���{/����Y�,Y���w�uW L7������6l�[��޽;~��Ĺs��y�/_?��O� �������>�� L9)��O>���<W��iS� ��T__���>�l�������>&&&�ޚ��r��M��P(�t$�P�B�=�PԦ�������8�W�������7�  �zHA�O>�D� �V�¼49�~��w��M  ����������ǹ�=�����2gΜ�`%��\YY әO� �"�S�6��Ç㷿�m? �G�o.m��V�z�  �mdd$���G����^7� �i-��|��Ǳw��ܶy���wܡ� �I�dɒ������Yگ��8t�P S_]]]<��39�^UU 3��;�7X�fM��G��믿�oB��H+�7nܘ/�,X  0�FGGs�i����  3M��:��?����裏���1֮]��v��;  ?X�}��������lꩧ�駟���� �I��E����������.�{ｼ%,�ݥ-�7oޜ/���X  0Y&&&�/�����7���"�uvv����cǎ9�~��w�1 ��J1`*�x���a�lfw�k4������=�\n�y��7��ٳ|��˗Ǐ~��ذaCno ����P{
u��  �ٕ������������sO,^�8  ��J�������Y�?��?������R�`
�?��Q]] 3��;�w�N�x�x��������o�>��GR�������  L����ػwo���� |����8}�t��Y݊+���"  ��m������?�{�7b�Ν>�� �r���?�y�b� ���;��TVV��w_����x��r+N___�l�Z����{,���  &C�ٳ'Z[[cxx8  �v���q�ȑ<i��U�V����n ��-[�,���/���ױm۶��H���J��=��3��#�D�P��ħV �`޼y���?�i\���C�iug�H7��b��Zxݺuy  �P��)mw|������u� 0	��>�;��϶��޸��[  ���*��_�"g%R!�R@��R�⮻�-[��w� ���;�$J!߇~8OWWWގ�w��]ttt�D�/��7jk `R�<y2>��hoo��1 �u��ϱS����}��ʡw  �.���ڵ+�x�hkk�ڥ������'?�I,Y�$ f;w�뤱�1�t>��q�������w�-�^]]]��jӦM�|��  ����ߟw�jmm����  ��ˋ�TWWǚ5kr�{�X  �V)��aÆ<iWƷ�z+>��S%�455œO>�?�x�c p��;�u��Z�n]�����sn!����������Aeee��*}q�}��&  ����F_|񅭋 ���������yZjsO�m�~��  �ŕ�Dwww�ر#�~���/Y�'�x"x��(
��I��@)$��xM��}�Q�ܹ3�=�����$������֞ښ���  &CjM�ϝ;�Z `�J�i)��}�����c��9x���  p�Ңɟ��'��3�䅔��=���\�٨��!6n��7o���� �L��&����[�I7	҅\
x���Y���S������O `2����ȷ��-��� ��#���>}:OMMM�^�:�X,  �Ej�N�i�����C^L�>7��,�ݿ����������o'�0466�m��������w
�sݥ�P�b���{�'���  &Kڱj�޽q�  `��E-����m�i��e˖  \��;��~���������������H�L�p��x��cӦM��� |7� SLڎ(mE�fxx8��S�{
���;L����JS{
�WUU  L����سgO�kk ��.]��w'}��7���2V�\�<�Vw  �YYYY�q�y����s��������|��9s������Q��
��O�`
K��+[t����]9r$>���܎s�ԩ�k������[sC{�J  \�� f����8|�p�[�;  �G]]]<��Sy�B��螚�O�80���)׳aÆ\4XQ!�	0|7�&R@���n����<����СC�����{�����?����ijkk  &��v  ��� �dhll���~:O[[[�ڵ+>��hoo�
�5�]wݕ��w�}�y �w�i���>�(�I7R���r�=5�\�x1�]�E�ڵk�"��*���9  �z�� �_�ǭ�>�`,_�<  �H;����~�O��A���}kkk����r��ӹ������: �~�f�����u[�l�x��/��{{{��%5�_	��cz  ד�v  ��+��۶m�� ��dɒ<���Ν�ݻw�'�|ǎ��0��{��-�h0]� pc��@_�?��S�����8q�D��I�S��CUUU���n��I�v�  �(�� �_muoii�͇.  ���y�O��<i����}
����/^��{o�իW� 7��;�,���M�N��t#!��Ӷ]'O�̏Ϝ9����͕��R�=mכ��[oͫ��B  �����w�ؑ�\'  0�R�f{{{���Q]]�=x��� �����œi�g�i��������?����_2gΜX�n]nh�뮻r���O�`�J�&���i��ӧO��4)�����/��mjjʫ�.]���)؞V��� �͒�v��n�  p�ŧ�~�}�Y��tÆ���  �}����r����/����{
�wuu�[EEE�Y�&��<+V���0	�pU:�O'�i�*m�B.W�Y������٩����i��4�-ʓ��͚���  ��mbb"��I��t�  7ZZ\�>~��s�}����Y5  |W�������I����ȑ#9�~��ᜃ`f+��p�J�=S���M��o���J[Ħ���I!�+��4.\������3+�
�EUccc477�c
�/X� �׬� `*Ja��;w������=  LiWѷ�z��N��<�]/ ����C=�'I��ʡ��G�ƩS�|V:ͥ���zk�Z�*�\V�\��^|��{K7�4��9ccc9�~%����J�nN\y�&�j�T>���������;�ܹscΜ9W�ijj�Gv  ��Ԍ�k׮���ٰ( ��itt48�;bnذ!�U  `���G}4O2<<���q�رxO� )��Ԕ�멝=گ���ϟ L� \7�B"5���9�~�&�䇆�b||���tA��U��k�&կ���ɍ�W�UUUy;������+�^ ��$�?�ݻ7o��έ `�H�2�"�_|1�ׯ_+V�  �l)+�v��<W�C:M��'N��ٳg���`)ױt���Ⱦdɒ���[n��0C����q%\~��x  �ۥ�v�ܙ��l� �t�v}뭷���2V�^�<�Hޑ  ���cX�fM�+R1ߙ3gr���Ǵý�����-�b�r�%�]�   f�tCe׮]����
  3���h8p <��.6l���  p#������R�=���?>O{{�������ei���������㦦�(++ f7w   �"5��޽;}ҍ  ���bδ���_�y��Ń>+V�  �R�}�ʕy�XZ��
I�����4�q
��݊Ҏ��]
�ϙ3'�9z:���tL��t�;wn �_"�   0ͥ#��=�W���  �F)��[oE�X�;�3���(
  SA
~�݇�|���n___�������ϡ����̏�1=ʏ��I�'###1666)������\���:�s��~z�����D]]]>���_�\O� ~(w   �i*x>����X��+ �����?�8>��X�fM�_�>**� `�+//ϭ�i�/_����|O�}&�%�_��W� {�g ���'9    ��ٳgc�Νy;[�v  ��R{��СC�hѢشiSn� ��L�: 3��;   �4q�ر�裏�ִ  ��I�iף�[�Fssslܸ1�ϟ    LM�    SX
��ݻ7>���  �����W^y%����G�e˖    S��;   �422���:ccc  L�K�.Eooo���Q]]�֭���?    ��   �����رcG?~<��  ����P|��Ǳo߾X�zunu/
   ��#�   0\�p!v���O�΍�  ��3::�;(�X�"6lؐ��   ���   n����������'  ��+�vSJ��/��7F}}}    p��   �ǎ������   ����R�]��_����x�Ǣ��9    ���   n��ƞ={��ŋ  Lm)����/��r466ƦM�b���   ��#�   p� ��������J����ƍc���   ��p   ��R�}׮]144  ����{{{㷿�m444�   \�    �lbb"����}�Y���  0��믿uuu�aÆX�lY    ��	�   L�+��O?�4FGG  ��R�{l۶-jjjb����jժ    ��p   ��R����>�������X   �K
���~��عsg<��ñz��    �p   ��R���?��;  ���P���{9�~�}�ŝw�    \;w   ��hdd$7�<x�jc{YYY   \��҂ؽ{��{
�   ���   �Q
�l߾=�9��  �&�:��?�����<�֭    ���;   ��Ha��ؾo߾���   �E
��ر#7��_�>V�^    �)w   �o���)|�F�  �CCC����Ǯ]���G�[n�%    ��    �g�}�w��-�   �-��}�ݼ[�ƍcɒ%   ��;   ��8p 7)��	  �����o��f�����?.   ��L�   ��/���;w���`   �H�.]�A��^{-cӦM���    ���;   0��8q"�o�}}}  p�uuu�+��MMM��}޼y   0��   �R[[[|����ӓ�  ��t�������ob���y�樫�   ��@�   �U�������}�   Lu��^�E��F����    ���  �Y���#��Qc;  0��k�3g�į~��X�ti<��Q,   `&p   f����x��w���-   ��tO�6���/cժU��c�E�P   ��D�   �������C|��� �%]�9r$Z[[��;�3    f
w   `�ٳgO�ݻ7��  f�t���Ƨ�~7n�+V   �t'�   ���}ǎ144   �E�z�w���.6o�---   0]	�   ���ӧ��ދ���   ��.]�����ꫯ�{
���;   �t#�   L[������o����  ��A����x�b�ҥ��OD�X   ��B�   �v���rc��'rx  ��K�Jmmm�����w�>�`
�    ���  �icbb"v����y~  �_���������z(n���    ���  �i��>�]�v���X   �݌���|�|�I<���x��    ���  �)�ȑ#�}��
   ~����x��ף��16o����   ��D�   ��.\�۶m����   `ruuu�o~�X�|ynt/�   0�   S���H����q���   ��:y�d��?�c�}��q���   ��&�   L{�쉏?�8���  �#]��ݻ7<�6m�e˖   ��"�   �t�O��w�y'  ��chh(�m������SOE]]]    �h�   �M��ߟ���Ν�K�.   7_ggg����bŊؼys
�    �Q�  �nbb"v�����l  ��ҵZkkk�򗿌����ڵk   �Fp   n��?�<v�����  �Ԗ�ݶo��~�insoii	   ��I�   �!.\�o��Vtww   �K��꫱hѢx��'�X,   �� �   \W###���Ɖ'��   LO��̙3�����w��ׯ   ��&�   \7{�쉏?�8���  ��abb"���G���{,�/_    �E�   �tmmm���.  ��ihh(�z�hll���z*���   ��p   &M
7���q���   `v��ꊗ^z)V�Z���B    |_�   ��سgO��U=   �˥K��ȑ#yG��<�-[    ߇�;   ������%���@   0�Ƕmۢ��9�l����   �]�   ����X�������   �U����u�ָ����{�   �k%�   |g��y�ر#��  �ϙ���={������'�����    �6�   �5����[�www ���(�]��,.Ey���𤋮����ңKQ(���2��~OMMM��}��先�?�ߚ�T�.]��|hh0.��/���h��\�M�cc1<2W�9���c� �����x��WcѢE9�^,   ���   �*�������-� 7B
�� z��cDMU1j�����*��������X�������ʊ�����b1��K�����beeT/?���,���4�QV������(��,��f�ti"�FF�>�A��O��������q������X����p������|�q�}�C�������qpp(.�fpx$�t�zKגgΜ��[���?k׮   �?G�   ���;��^��� |_��2�����p9�^S,Ɯ9�QW[uu�cMm���Du���zu�Kϋ��L�Sz^(��l������W|��dI�F��r ~xx$7��c鵡��.�P����?0�}��S������o |ccc�}��طo_lٲ%���   ��  �?��ŋ��o���� ��Ԭ^,/��,*J�k�����>�룮�&���Ŝ�ڨ)=����buMT��U�c��:7�s�
��.�{J�]������P^,�;���`i��b�_����x1zK_��틾�{�@���/��R�Z�*{���    q�    �{��ɓ]�}�eQ����XQ�ڪb4��ż��Q?gN�ח�nN���Eu����%-R�-��H3����?>1C�����w9��ן���7:�����?�zz�b�= �|i�ӑ#G��ɓ��OĲe�   @�   ���ٳ��[o��U f�BYD��<������be4ϛ��^���������S��)�\QY��򨫛�g�_x���H���F�Ł��닞��|����=�q��+�GF��a��}۶m���[�l����    f/w    ���r��ĉ��V^V��<5�Q_SM�Rp}^�K����������!���(+�����X��������DoOO���EWww\(M�����s��14< L/����[�n�x ���    f'w   ��Z[[�wމ�Q-� �EE�J��<���PW-�͹����1�4̍چ����vf����<-��_����N�����t���������	 ������裏�������F}}}    ���;   �Ri������ L-eeeQU��W����ǂbol����b�ܹ1�a^�WVU�uUUձpѢ<lhh0߻.tEǅ�����;�t��� n����x饗��;����   0{�  �,���o�ccc�͓zի*ʣ����幕}������%�����)7��k�U5�L���X�(͟���GggG�?��:���s��8���.]
 n��}w߾}q�رx�駣��)   ��O�   f����x��7�ܹsZ 7P��,��s������X�2?̟s���~^c4�+�P(��)VU��%K�|U
�w]茎��8{�|�>{.N�k����w^p]��/��W���{�t�T   `�p  �Y�O>��>�(����룼P��QWY5��+VDKsS,X� �5��ܦ�h(M]}}��	f�t���/�s�W^����=5����S9�~.�/��;��:r�H���ŏ~��X�xq    3��;   �p�����oDggg 0y*R���<�)VDS}],Y�(���4�DCSS���f�bUu,]�2��J�.��F���ўB���ƉSg�����{�!����5�ҥK㩧���   3�;+   0��ٳ'���D ��e9�>�X���X��%ZZ�������9j��@RV�5�an�[V������pt�?gϵ��3g�ę�q��#F���%�w�k��g�&��>�x�X�lY    3��;   �@]]]���G___ p�
eeQ]Q�f�,����X���Fc˂<��GyEe |W�UU�xي<|����htu���z?{6�N��ֳ�h4ƅ������ضm[,X� �~��(�   L�   0�|����'�h�)�^[Y����^U��2�9���7�,��M�R��~����EK��u�����;ݝq�T[�:s6ZO��g����� �����غuklذ!V�^   ��&�   3D����o���@ 𧊅�h���2�^����/\��_ifof��B��ۤ���˯ƅ�sq�̙hm;�J�����@���X��������3�<UUU   LO�   0ͥ��w�y'�;���K�B�I��U�cE4��Ăŋ�y�hZ�8�,��� �.����+n��ࣗ_����Ϟ��S��h�8q�\����D �V���������o�=   ��G�   ����������P �V兲��,�9iR;{�����/�����ļ��(+��I�����u�x����h�\舳�ڢ�d[n=�}�d<&,�f��������������Fuuu    Ӈ�;   LS۷o�}���l�����1��27�ϫM��K�)��/X�[�+�U0�TTV��.�s׃ǥү����8w&�N���'�TGg���؄�;0�uuu�/�7n�U�V   0=�  �4�nп��kq��� ����hHa�bE��sr�}��%_��/�B� |]ڹbn��<��'~Tzmhp :Μ�S�Nű�q�ԙ���q�w`f���{/��?���Q,   ���  `����O>�K�������<7�7�c^Ue�k��2̞Z��ļ���໫���e�n���Ãq��\�=}*�;G�NG��h���L���[�n�'�x"V�X   ��%�   �@������ 3͜b��v��U����e�}i�,^����QUS�Wޚ灍���{Ǚ�q�T[o='Ξ�����8:a�%0�6���~;�-[O=��]�   `�p  �).5��ڵ+&&&`&�/Vļ���[]����0wn,X�<O��e�]��#ޗ�Z�g�C�q�T[�i;G�����=2���������矏'�|2/^   ��"�   S���@�������� �Ϊ+�s�=Oue���F��e�p��XP�����Ԕ-_�6�#OF\�뉎3g�ܙSq���8}�;��Fcx�bL`z�7�x#V�X�7o��   S��;   LA��۷������BYngO���h����%KsC{
��76EY� �OZ��f��u���~=���v2N�8_k���C�72��`��t�R���Ư~��زeK455   p�	�  ���^��8w�\��0�ʢ�x��}^Ue4��y��h_�tY4-Xee1f��Xi^sK���=O��EǙ�q���8z�X����ޑ���q��688/��r�~��aÆ    n.w   �">����v`�+��E}UE��2Ԟϩo��V����ce�* �]��+�π4�=�9����q��X9v4��^������(�v�ԩx��g���>   ��C�   n����ضm[�8qBk;0eUʢ15�����TUV��ũ�}EnjolY �U�5��r�</MDwGG��:'����'�kh4���bd|" �����x饗��{���?   �O�   n��'O�[o����0����E]e!������U�Q����E�WFEe1 �Z���b�4���P���q��h=z,:�rؽw�nF�͗��ݻ7�;?��O���6   �G�   n��������_|���2*
e����4M���*��e+r�=Mm}C �d���������x��j�3�����cq��B\����p��<�����/ģ�>k׮   ��p  ����;^}�ոx�b �l����\S��U1��2�kkr�}��[��pC
�WS=���q��'���9��#�32�#�p���۷o��Ǐǖ-[J߳
   \_�   p�۷/v�ؑo���ee�PU�[���������@����b^KK��~��RW?7��}�G����8}�H?v,.E��Xt��rw�F:s�L��?�c�ϟ??   ��G�   n�h����ԩSq�$pcU�rK{
����ʊʘ�xq�/�uM���	 ����kb��uy����q��X�;g�z�sh4���b�96p�+��w�yg<���   \�   p��;w.��Ӎp�%5�7�TFSM1�UWFuuM��Y�lETTV L'��W�=�ēq���8}�h����sp4:��bd�nI�����hkk��{.���   �\�   pm߾=�������幩���"�VUFM]],�eu,�uu�,Yee� �� �L[�ty��6m�������#q*��ϵ�f����v .�  ��IDAT������կ~�6m�[n�%   ��#�   ����@޶���' �������,�P��Ҥ�{��h_��X�d�P; 3^Y�Wc˂<w=�1.��ę�c�v�p�8y2������`2���Ż�Ǐ�͛7G���   &��;   L�Ç�{����p=4TU�@{K]UeQW�KnY�V�M� �Vu�sc�����j����S�98]C��3<�X&Kkkklݺ5�}��hll   ��p  �I211۶m�7�&S�,����5��T��B!�6��M��V����� &���H\����xi"�FF�����t���/�����<^��x��cc��mtx�k�/�~��|��+�7)��GEŵ}��vq��,���ߓ~oR����g����/�^Q,�]"���+K�w**��+K���ǅ���π��a����h;�Ei�����04�����d��_~9x����{   ���  `ttt�k���ohL��Ծ��*Zj�Q^(����X�zmin�9s��R}���xdd8FGFJ3c�#9t�B�iF���|<r��ޛ�c�D��+/��BEy�U��9_���)9_����=�yeUuا���b�ZX�"��\���y�{{.�ݏ|���5<v��]���.]��w���S�{�X   �p  �h׮]�w��|#��Hm����_S�uUQY(�a�h_�f��vf��A���H��xh����/�P���3.ޫ.�߿r����TU�DUMm�X���t,��ǜ������yz�.��#����Cq��+�h�������[�n���z*�,Y   �w#�   ����H���q��� �!j+�cAm1Ω�b�,j���@{jkolY0SLL����`ib(����p�8<4�/�K����.)$�f���OZ�B�Ś�|��������{u
�פ�5QS[�)�?���)�Z�!υ��rн�ȡ���C�����266o��F�\�2�|��    ���;   |i���~;߰�>R����X����(���Ukr��y��(+���bbb"�.�������+K�����_̡�^O�0��"��/L\��򊨙3'�k뢦�.k��DUm�׎�����Բ0Ͻ��3���������1�;Gcpl" �U����^�����Q[�9   |;w   ���o�����*|gU�XPW�QSQ����޺:��,Yee���&��^�X��+=���)Ȟ����S㺟�L��c��ӝ�/�,�nW��W��7D]CC>
��li�Y��yx�Gq��8q�`�>v4���s����h��߮�t���/��͛cŊ   �e�   p�FFF��_���� �V�BY����9Ŋ(
�p��X�v],^ykn��)~SX�b_OiJ��t�-��{��f���y��ȅ�����I;o��{m}×���W�5u���=3C�P�f���#_D�r�{ϗ����؄�>�7�;��\�2�|��    ���g   pN�>o��F�����)��ESMe,����ұ��ZCSs��m]������itx8�sp�4����@�qOOne׾�]Z������?���Kǜz��C��q�c}Cng���,�-��ʓv�8u�p;�?�:�G��x��ą���m�&�����K/�s�=U��   ��p  �o�}��ؿ�����cAmUnl�,�EMݜ�Ծ�u���p�\�4�ep�;������+�z�s� ;�iaI���<,�ޑC�s�E��ƨO��ω�yM9���~ί���<Ο����Ç���@t�������?�[:oۺuk��G?��˗   �u�   �R[�?��?������T�r�}aij*
��u٪5��ۣe�2�L����ׯ��{R��+�'&&���Ǣ��B�?VUS�E͙�)�^z\?o���)��ea�{7>gO��C�Ǚұh$�ӌ��>�����x뭷bݺu�裏   �/�  ��hoo��^{-FFF���ʢ��2�V�cY�����s[��[WGyEe��511�C�}]]��}��0{O��t���h 3���`�<�O��������˶�yM�ϻ<�kL�B!�ܲ*���@�8|(��=:�{x,�/�f����8�O�����U��    �  �O�޽;�����N��H!��bynjo�-Fy�yjӽ��;Jsg�Ω�.R�=��s�sg>� djc�3�c�����|��J?�jJ?�����mj�y�[r|�P�<U5�q�=���:�������Pt|���;< ����u��زeK,\�0   `����݇wTס����M�����@�M��N��o��%\�Yy�ɻlc�m c�cS%��*H��4}Fq�QT�|?���b��،�>���&�    �7
��z{{599) x��4����v�Ô�phs[��־iK���S��/��>�^���� ��� &_�����[�wk�UM4�H}�"u��QB������^��{�ɑ{Jds�N<
�g��^�\N��v�ڥ_��W    ��p    �hffF~���� �4E}.m
x���jcuڶc��tu���
�!�Ĳ�g5,/���!����� ֝���_����з�{|>��?�jc����ُC�m����sniﲇ�(a��n]�B[B-d�Jd�0�?5��d}v߸q�^x�ꫯ��v    �jD�    P���ǟ�9�C v[��Ծ)��4�r��ұ][�w*��$ౕ��K�Z��f�5��Ѱ� P��ɤ��F�����DU��-�Vۻ�6������h��~c7�[����=2�+z��hr9�4��@U����;Ｃ?��Ojhh     Ն�;    �j
?~\���ہ*��m�Vȯ��Y�v�Rs{�N�U�\6���3���������̞�� ��:^,~�YC��~�
�[A�hCc�Ѿg��g��[��ܦ��G�nZ݁*�-�~��G��/~��{�
    �j��9    @U���Woo��� T'�ӴC�߶�{<�ڽK��(T�S>������4�`�ne_Z�g!��d�J11<d�ǂ5��44*Z�h߇c�r�\³ki�ԍ������Vw��YǠW�\����x���)     �w    @չy�>��s��@u��v��L۾s�Z;�	�U�������v�}~fھ�`J�|^ ����`��;��s+��D����ZM�ֽi:�'
GT�=j�����mvvV�����^{M�pX     T:�    ��r�����@u��v�é��Nu����<��_���ķavk��9 ���.l��1��~�j�#�56�n�f;��Ddo�aV��͟�?F�;P��鴎=����C     T2�    ����d��sssPC���`{�����hL���m�9]n�r��	�NNhvjB���P{.� `�Y;%=�ݺn���x�oP�q�bMM�54�s�hi���K��k�mu/��TN��i���Zt �2Y���}������;     ���;    ����̨�����|VC���nۭ�v����vm۵[ͭ��V�������v#���};��{H� JH6���ب=,Vy(��彾i���U��⟅5�?���ud�:��4���T"�\���@���u���kr�Y�    �<�    ����:{�,!G�
]5��j�e�|��:��Ӷ�����ʑͤ5;5���1;eڧ�˲�	 ʉu|��-�P��6ہ�ئ&; _M����O���߼Sm5^���$3�XJ+�+@�v�{��w�{$     ���;    �b�9sF���P�b>���E�.�y]S�:��S��)���f����� *�r|������n���?�Ge�U������?fR��m��LN��&�PY���;��������     ���;    ��Xx�=j���L.�Ц���{��Z;��s�
���R�Y���531nߧ�	 �O&����=,�áh}�wB�V�R�F�
G�_�yL��i�TMAS�M%2�X(T�B�`�\7==�    �J@�    PQfff���k��T��ˡ��W~�LÐ��W���صW��c�������F5U&ƔN& �+�󚙼o�>]�_�j�вE�-�jl�"�ǣr��ީ[W.����:L��x�Z<�z��hb)�D�  �a``�>'��k���v    �rF�    P1nݺ�s��ie�6B����)�Q��_��7�s�~���4M�|�������};�>=>j7� �,���u�F�!\W���V5���-��./夥�k��c�F�����&�3�Mf��Y;ٽ��v�=�    �rU^g�     �gΜQ� T�i�)�-��S�á֎.;�n�Q�@���=Ӄ�q�L�W.�. ��g-t�{0m�����p{lS��7����EцFFi/����)X������_��i�T���匦��
,ʙ���ѣGu��uvv
    �rD�    P�_��Z� T��a�ڭa��.���إ�/�(_ (�������Fih l�|>g��ƍ�*S�kܤ��-�k�\�����N���Һ���ijk�W[j��Jdt)�t��;P��?gϞ����t    ��p    ��������!w �/�v�9�S��m?��jԱk��w���JW:���٧�P���E Pjr��7?�F���"�Xc�xohnU��^F��Z:��=���Y��o
���x<�0���RZKټ �������k��&��-     �w    @Y�u�Ν;g��(_�a(�u�9�Q��e��kP����ҵ�$[U!�sY�LM�-�V+���>� e'��|'����T�Ԣ��m�\.��,����kia^�x����e��LN��2v�@��v�{��w�{$     倀;    ��9sF���P�L�P�߭-5^��;�n�ɶ���Ꚛ�Ҳ�R�܃i; 8=>�٩I� *K:�����=�Ex����ukq��{�{��]��RP�v�&�T"W��g��(/��wG�Ձ���)     Jw    @��f�:r���7����q���n����.>6�vt�{��T�
�#�J���1;�>1<�TbY  Tkg���	{ܸx^�O��[��ҪM[�������w�L��1��TWا-!�&�3�Jd�+uʅ��v��Y����7���     (e�    e!����T*% ���0���WNӐ��U��Աk�<>���V����)M�kr����n�`  ���_�������ݭ�{��������g5�B5Z�/��X�um5^���Y��S�t�F__�r�7d����    �j!�    (y���:~����� ���۩�W�~���s�ϯ��{յw�\n���2锦�Gii �)X���`ָu墜.��m۪���[s{�����Re���p����l*��xZ�s6�������ӡC���0/    ��    ��v��5}���e&�q��Ƨ��e?�#�~�EmپC��6-�  ��\6k/���6Vg��7�mS�q�3���tt�t��1�0T�s�����tN�񴖲݁R����w�yG�������    @)!�    (YgΜQ� ���ץ�Z�B�G���u����K;�e��XoV�njlD��jr�ҩ�  ��Y���G�����|jڲ��7�l��ޟT��A�P��E��0+Zc1���bZ�{ �+����?��~�;utt    �RA�    Pr
��>�����@y���j��~l�۴��oj�J�}��	M���M�VS�r  �/�L�^�M{8N�55�a��m���?���1T�|���MM�pw����_��a�c�TY;:}��g�9��_~Y     ��    ���H$������ J�������֧��a���Ҫ]���b�M��Z�/؁���w4;5aU  @���s���ճgT��i�Vm�ڮh�\���Y��Ǭ�{Mԩx&��4Aw��ݾ}[�ӟ�$�4    �F"�    (����裏�-��.+���V��尟�tti��_�6V'�����f&����A{,�  ����Y{�]�,�F�۶�i�6�7�|.���V�{ryI�,�vhGԯD���xJ�I��@)�����Çu��!��n    �Q�    JB__�Ξ=�B�  ��0�z�G[j��9�[;�k�/)�k/��jr��h�V&�  (����\��.�[�Z۴yk�}o��_��J�w�����F��� ����%���;z�7�    �F �    �p�}��p_YY��c��������B���Z6������hjtD�<�\  Pɲ��F���jr�C�4Vн+�Skȣ�xZӉ���#����ѣz�W�u�V    ���    6���~��q���	@�q���n����v�v��y[�v����k,�N�j��؈
��  @���LK��T��1fGا�G�iM.tJ�����'�h~~^���     뉀;    `C$�I9r���@i��훃^;h�"ؾn2�&��j  U��4���W<�hl�Fw��@I�ꫯ4;;�?��    `�p    ����رc�d2P:L�P�߭�Z��K:�����P��ݒ  P�<V�{�X��
�ǿ	��F�v�{����׿�UN'    ��c�	    XW������O�BP2C��{�V��3M�Ԗ�;���_+�VWryIc�w4^�S|  �;��w��L2�1����;���7�T(     k��;    `�\�r� J���󹴵�/��ߍ�{^����aa�d�i����'G��  x�1jWا�G��f�Y�8���jr�ӟ����&    �V�    �ũS�488( �!�s��֧��a?oli�����±zau��9M��j�������   O��4��+�i|)��)���F)
:y����G۶m     k��;    `MY>�?���1�x����S��贐l�����o�_�������>>tW�,�+  ��*��:���i4��B:' ��:�s����q�۷O     �6�    �5��dt��-,,�ƪ�����Zϣ�A�MM����75�g�x{85����ӧt2)   ���S�cNͧs^Li9�N9�F���/�s>���     XM�    kbiiI���R�� l��rK�OQ��~mh��~���-�󙝚���~��P*�   �W��T�>���tO*�+������/�i�    `5p    �������(��
���j���ﶟ�D��������)�xóI./id�OC�ohia^   �x�SaOPS9��SJt�����>�������I    ���]    V��ȈN�<�B�@�<S[j}j��e��5����ߪ���`�3�e3�;�{��5;y_+++  @i��}c>��^�������䙗�eaaA���:$��/     �w    ���q�>��s�p��ZB^5�|*>���U��_�k�~��Cx:+��éI�뻥�;}ʱ#  @Y0����b�:�K�����i噣�"�J����z����F    ��"�    X�Νӭ[����Q�ǣ��>��N�:������\n��t�jlp��'�  @yr������\v��T"# k/�˩��G�����,     �w    �s�׿����AX_u~�l�92C[������ˤS����ۚ��/   T��TGا�A�F�i�&ٙXk�BA���?���/���[     <-�    �gf]�<r�fgg`��x��V��-�������[�?)��krdHC�ojjt�~  ��e-
�����ix1��l^ ֎�������E��׿     O��;    ���R)���{J$�>�.��j|vs�%ڰI{�;�7����ZZ��ȝ>ݺ���   P]j=N��M���R9:k�֭[������      �w    �S�.L>|X�tZ�a��r9L����\�߸P8�ݿ����;���;�s���&��4t뺦���&A   T��ϥ�ש�DV#�)�9F���ؘzzz����4M    �s�    ����z{{�ϳ�;�����A�Zk�r|��$�Ш���d�~��̴�nߴ۳�   ��d���n��\_J�~qs����]�p��!��n    �S�    ��ݻwu��i
l��%+ʾ)�Q[�_.���v�!�������h��u�=�   �s��c��n��}&��շ�����{O����+��/     ~w    ��u�Ξ=��m�T�ǩ�H@��{���r���K�>+�n��G��)�%�  ���u���ks �������\��L&���_o���jkk    �!�    �YW�\��˗`�x����j���V�-�]r�����l:�{}7�`{|~N   �j��[�L*�{Ie,�VS.�ӱc��ꫯ���^     �7�    ��t��y]�~] ֆ�0�R�UK�'���_�u�.��v   �=�x�^�s)�uj,���rFv4VM>��G}�����jmm     ���;    �G�>}Zw����������?'�(��I�*��ibxH׮jvrB   �z����x��wih!��tN V��ʊ}�������     �p    ���ǏkxxX V_��T{دZϓ���ڽK�U���yݾ��[7�I�   l�ӡ]��p����\^ ��r?{����v�b�2    �#�    �Q(t��1MMM	��r�������>��F�뺺U-VV
�֝�W5=>f   �R�8��>��DF#���U��p��%�R)���    ��;    �[V�������ܜ ��w�1���Z�\󩿾�m�|��*]*����ۺ{�k%��   J�Q<�o
�U�sid1��d�E��*�~��������V    ��F�    `�f�z�w���$ �'�q�=�W��x�ﱵ���i�{0m����  @�p��:�>m
�5��T<���300`7�<xP    ��E�    �d2�w�}׾�:|N���^�w?�����ڴe�*M����{���K�NM
   (W�bֽuA=Hf5��R&_�g7::�?�P����     Չ�;    T�x<�Ç�[@x~�!��������ںw�4MU�T2��[vc{ryY   @�����85Oib9# ����:z���|�͊�    �w    �b������Q.���W�q�3���X��ٶ}�*��̴�޼��������  @er���������|RKټ <���99rD���I�    �	�@    �Rccc���U(�u:��S푀��U���MM��DU�V����{v[��ب   �j�w��[ЃdVË)e+���<��[o��^�97    �tp   �*t��]�>}�p;��Ц�G�a��Ըڶu�R9�f����Tb).   �Z��\
{���� ����L&��_��W    *w    �2�n��ٳg��B{�<Bn�:#�<ksz��r��c��I|a�����V>�    �e�������bJ��́��N�u�����
��    T6�    PE���k]�pA ���4�V�SsȻ�����e����܃iݹ~U#},�   ~D�ǩꂚLd4O���3�Tr��zzz���+�
    P��   @��z��.^�( �.�s�+��a��{m۱[�l�x����W/ivrB    ~�aHM��V��BJ�iv>�F>�Woo�^{�5���	    P��   @�r�= <�ˡ�H@��4���E7�
y����//*>?'    O��0�3��\*��Ť�y�܁'U(��G����    �<�   ��}���ꫯ�陆��oq�����jo7�~��$�Ʉ�޼��׿V:�   ���:U�j|9��Kis��r?q����?���I    ��B�    *؅���_�ӳ��;����u}_�0���[�biqAw���[ו��   `u9�� �Q����bJK�� �<+�~��I<xP---    T�    P�Ο?��ׯ��q����}j
z7���ڶ��h��NM���eMie�I   `�\��5����bJÁ�e�WO�:�����jmm    �2p   �
�駟���O �N��VW4 ��ܰ�ö����`��//��v    ���ѩ��V����BR�ivQ~�r?}������jkk    ��p   �
��'����_ ���4������߇��Wc��_�_)�&���֕/�pzJ    6��ahgԯߴ��s~�r?s�8���    �w    � 'O������Ө�[��A;��ںw�4ׯ=�
�����K�8�P    JK�ϥZ�CC�)=L���+�~��Y�1!w    (o�   �B�8qB����'�q��*�u�Tl�޵.�S(�5zg�nl_Z�   ���.�]�#~�&����Y�Ν+�{���    �<p   �
p��q��i
z���al|k�cu�6+���{�Y�뻡����\^   �����=N��ӚJd��YM��ϟW.��Ν;    (?�   �����j||\ ~���PW$�p	��?�u�ڵ�g�)ݹ���\��~   �<9MC�^E�N.$������K�.�a�]��g�4    ��!�    e�p;�d������j}2K���1�˭����:=�L�m�C�����    *C���uA�.�5���!^ �e���B���|��^    �|p   �2T(t��QMOO�O�ꎅt;T�Z;��t�^�|:�P��_ڭ��\N    *��4��ƫ�ץ�I%s��������߿_    ��@�    ʌn�������q�!��������l���;Vg�t��   @�	��W��RF����]V��ڵk�9�_|Q    ��G�    ʈu!������� ���۩�h@Aw���#�6nz��A�   �n�a�-�Q����\R�<m���B�ׯ_�i�4�   @(���     ���v������ڭ���Z��(�v�.�����J�   �
�z�>�1��}9c�z����n�^x�    Jw    (���z��� �0�ӡ�j=.�����O�u�   �k��87r��|Ri�܁oY�>���k{>�o�>    Jw    (===�������=��,����6om����_O�   ���u;��.��xZS�� <b�ܯ^�*�ө]�v	    Pz�   @�����߿/ ��u:��̈́�hk��]H�������ו�l   �d����Z��V��BR� <r��e���;�~g5    ��*ϫ�    P%N�<���q��:�[ۣA;�Q����M[�~���Yݽ�n]�X|L�"   �g�:r5����TV 5����cB�    PZ�   @���?����!�.�i�+���l�]2��Y>����v�=�L
    ��5���4�tjp1E�;���/��r���C    ��@�    Jп��/
�w��=���r�*wm�w~�B��ᾛ�y�����   ���t;uw>��LN@����Ϟ=+�0���.    ��#�    %��O?�ݻw�ߜ��ma���^U���f�o��o�wt��9--.    ֒�ahW̯�DF�S���r7MS[�n    `cp   �b]H�����x]��S��m۱˾�����t��y-��    �S�߭�ǩ���♼�jf5�[�N�S---    l�    P"Ν;�[�n�� H��5xد͡�hm��r�y[���G�����   ��b-&�hl)��xZ@5��˝:uJ$�    ��;    ���/�ƍ����Ю��.�*M(�g~���q   @)0��5�Q��T�\R�|A@��B�O�֟��g566
    ���   ��t钮^�* �4<��0U"�   ���ˡ}u-�4��
�V�BAǏ�_��544    ���   ��ꫯ��p9Lm��    �N�PWا�ǩ���
+�����8�^__/    ��!�    �
�_�xѾXT�Z�S;�Br;L    6^��e7��'����FV�����_]�XL    ��A�    6��k���_�vFql��iK�O�a    P:|NS{c�/�5��a�>����o��p8,    ��#�    �l``@.\P�<�nm��pz    J���%�����'�)rG���r����[o��`0(    ���
2    ����}��'4��������i�    ���ǩꃺ3��\:'����y;vLo���<�     k��;    ����I�8q�p;���4�	�!��`    (7��nGԯ�匆S��M&�ё#G����Mn�[    ��A�    ���̌z{{U(T��ǩѠ|.�     �)����Jd��I*�ROO��z�-��L    k��;    ����e{�bkc�����W[�~    T��Ԟ�_��)M'��I<�C�    `�p   �5d5:���{�f�Ћ��r��*�u	    PY���Z�"��.$�+��sss:~��^}�U    Vw    X#�LF���r�Q�ǩu!yl�    �,�u���>�D��P=&''u��)<xP    ��C�    �@�P��Ç�H$T��W��C    �*�s��hh1��;١z����ܹs:p��     ���;    �������E��i����    �����������BJ����Ν;�x<��/)    ��#�    ����W>Pm�n�vՅ�u:    �^�>��.���J�
��͛7���={    x>�   `?~\�MSЫ��_�a     ���޺��Χ4��
�t+++�r��~����    xv�   `��={V������0��!�     �ɚ3n��4�p��bZ�����>���VKK�     φ�;    ��˗/�����thw}H~�C     ��F�[A�S}s	�������z��W���     ��#�    ��ƍ���/T���jn���     �9��}u�]H�a*'��
�8qBo�����     O��;    <����?^+l��*aRg$�MA�     x�⤲;���rF��8��J�����ӣ��zK�`P    �'G�    ���ȈΜ9C�U��rhg,����	    �g�p+P�c�%�)p^��q���ߖ��    ��pE    ���̌N�<io7T��ϥ��ݶ    ��q;�B}P�sI-dr*U:��|�����2MS    ��G�    �R"�бc��&�������'� �    X=�"�1�F�i�/�T*�|���~��!    ~w    x
�\N�V6�P����hPu~��    �k)���G~���)VVT���9�:uJ    �p   �'T(�p�ոT:�ˡ��!��    ���|���T�\R�|A@%Յ���/    ���   ���������J���[�    �^.����?��B&'�������F;w�    ��p   �'p��MLL�t�5>m���0�    ֟��zg̯�xZ�Ki�feeE�.]R Ж-[    �>�    �3�\����>��a�U�w    ��d-�����4uw!��ʊ�Jb�ܭB��^{Muuu    |w    �	w�ܱ�@%��]���     ����*�UM��%��T�B���Ǐ뭷޲��    �F�    ~���>���Q	�T1�[ݱ��<     �&�rh_]@�sI-dr*I.�ӱc����o��fW=    x��;    ����E����MJ@�j��ik�O�A�    P��E�;c~���_J�$�tZ===v��i�    p   ���d2z������T"�i�;T��f0    @y��fo	y�w�\H)ώ{� �x\'N��_��    �   �wX�����ݜT"�ˡ��5�9i    ��:�˞�ޞK*�g�=T���)}��z�W    Վ�;    ��#G�؍I@%�x]�Y���    e,�rh_]@�&��e>T���!�B!�߿_    P��   �7>��#����DMA�:#�     ({.���X@�I=HfT�k׮)���S    P��   @����5::*�uDjy    @%1�3��ij4�P	VVVt��9;�i�&   @5"�   ��Y�Hׯ_Pi����!E�.    P�Z�����̧TXYP	N�<���zK�PH    Pm�   �jccc�pႀJ�s:��!d�    P�b^�<1S�&�-rG�+
����?��9�D;    TfA    �V<׉'�m�JR�qiW]P.�)     �E���޺���Z����L&�cǎ�o��    ��p   P�r���9b��dSЫΈ_�a    �j�q���B�	ͥ9�򷸸�S�N����   �jA�   @U����L&T��Z_q�    @53iGԯ�xZ�Ki�nllLW�^����    Հ�;   ��s��	���
��Pw4�:�[     ��-!��NSC)VV������׮]SMM����    ���;   ��b5ݻwO@�p[[�ׇr3�    �5�\��η����|Y!��g�*+�
    *W�   T���!]�tI@��B�V��
�    �r;��.���J��ʕr�裏����]^�W    P��   �
sss:u�}��~��cA��     ���:L���7��b��;�W.�SOO��~�m�&�    *w    /����ѣ��x����=�A�    �'�4��uw!��dV@�Z^^�ɓ'�ꫯ
    *w    �P(�ȑ#J��*���_�5>    ��g���>���F�/B�����_|��^zI    Pi�   �h������;�|w,�z�G     ���=r���ZP�n߾�h4���N   @%!�   �b]�xQcccʝ������z��    �Z�.{�}g>��
1w����ϫ��V���   �J��q    ��ݻ�ꫯ�;��Ԟ��]    ���:�+�׭��rB�(?+++:~���~�m��~   @% �   �������������\�m���a
     ����8����Ä����r���u��1����ir	   @�#�   ���R)����P�b$�[��Ү���!     ���S�c��%��������_]    P��   �V������d2�Yc���Ѡ��     ��ihgį����R9����:{��~���	    �w    ���WKKK�Yk�O��~    ��g�#���BJS	JP~U__��۷    �w    ���˚��ٻ�/����㯻�]f�aeSDC�|�6mOlN�tM��&��6�Q������ *"3,�,�ܹ��&]�����<�|��0?���~���ʕ@7{tC_��   ���C����\�=�&�V+'N��ƍ�iӦ   t#�;  ��>����W�
t��:��M�X�	   ���UR.$ߞN������^�O~�T*�   t�;  �����s����C�F�R1On�@�+:   t�ͽ��|���������Di4���~���~:   ���9  е��f����m���Q�\ʁ-��W�   �i�ZΓ#}936�FS�N�h��=z4O=�T   ���  �Z�=�\&''ݨ^.��[S-��  �����v�>:��;]�ټys��   t�;  Е�z�\�r%Ѝ�+��<0�9   ��7�}mS;r���\3�-N�<�M�6�?   �@�  t��>�,��կ�h�֓'7�T,   �.��ڑ�ٱ�L���A��ʡC���3Ϥ\��   �ϛ  �U�����/��@��W��@��   нz�z�bco޿1���;�avv6?��O���O  ��	� ���l6�a�F��l�汑�h�  �����<9җnLelz6���!ǎ�w��   t2�;  �5�{�LLL�̓�����+n  �5����؆z>��|9%r�;�?>�6m��?  �N%p  ��[o��+W��͎�zv�   X{ڑ���zz��|>q7�N�<9��  �N$p  :�g�}�_��W�n�gC_�   X���\L>���Z�V:�g�y&�l  �<�T  ��6>>�_|q���E�P�c����   `}x���R�����}ˢ����������/��/  �4w  �c5�����?M��t�R�������^	   ��<�ۓr!���T$�t�۷o�رc��w�  �N"p  :�s�=����@�(�yrS�j=   ֧M�����|pc*MK�t����g���ٷo_   :��  �Ho��V�\��=�b��e0}=�    �ۆj9�o����ij��p���/�#��7  �� ��s�ҥ��W�
t��b!_�< n   ��P��'6����̩��`�V+�3�<�rYF  �>o&  @G���ɋ/�8�ݠ����^q;   �TJyrcoΌM�!r������СC����   �6�;  �Q����m�0�A��q{]�   ����o���c�����������5���o  `5	� ��q���ܸq#�j�RlH�,n   ~��_G���t��n|��lݺ5   �E�  t�O>�$�Νt��,����    ܋����FzszԒ;��^�O~�T*�   ��;  �ꦦ�r���Z��|���?�:�JI�   ܟ�w�'G���g暁N�h4r�����?�s   V��  Xu?��O�M�����r`��   X�z��'6����d���P7n�ȉ'��o;   +M�  ���_~9�n�
t�v��uq;   �ڑ��#�9=*r�s�;w.=�P�o�  ��$p  V�G}��?�8���+��<�q;   �D��v�ޗ3c�n���LG�ɏ���j�   ��;  �*����ꫯ��j:Y��[�S,   `)UK�<��7g�&3%r���������я~  ��"p  V\����~�����d���r�`J�v   `�T~��>:�I�;�֭[y�������  X	w  `Ž�����Ɇj=��恔
�v   `y�o�{b�/g�&31k����f۶mٹsg   ���  XQ|�A>��@'����M�v   `��G�{sF�N�:v�X�lْ���   ,'�;  �bnܸ��G�:�`��'-�   �������щL5��N�l6�����_��_  ���  ��h~<��s�?�ST�9�yP�   ��v���H_N���@w�ܙ1yꩧ  �\�  ��8x�`&''����oL�(n   VW�ȝv�<��Cٽ{w   ���  Xv�O�ΥK�����4����   @�hG�O����wrw��$���Z6oޜ���   ,5�;  �������o:UoO)_�:4h   �I*�K���K�w�,��9������?��O  ���  ��ir<����?��˥|}ˠ�   �X�R!Ol읏�g�������9v�X���  `)	� �es���LLL:Q��?��J�   �NV+�䦾�w}"�"w:����cǎ<��#  X*w  `Y�6.^��D�C�v�^�   ]�V*�ɑ��%w�;����m۶T*�   ,�;  �䦧�s�ȑ�Z��<���[���   @ש��ٿ�7g�&E�t���������~  �� p  �ܿ�����h:�|ܾup~�   �����#�3c�i���cccy���o|#   �%p  ��ɓ's�ƍ@��)���z�   �n��#�9�;��w�͎;222  ���  K����9u�T�������-�v   `��oG�zs���D�W��ʳ�>�b��  ��	� �%�l6���|�:I;n�������  ��e�R���#ro�.G���ɑ#G�W�W  X(�;  �$���LOO:I�Xȓ��W��   �M����G'"q�|��g��㏳gϞ   ,�~  `����\�|9�I��B��4���W_   `m���w���nM�a�����g۶m���  ��r�  ,ʝ;w��k�:;��l��   `=�T��\���ܲ��k6�9t�P~��  �~	� �E���~����@'yl�?�{�   XO��V2;��gw�Vۭ[��_�"��  ��!p  ��ѣ�}�v����З���   ���}�:�����L`��;w.;w�̖-[  p��  ��|���y������z��   ��=2XK��ʵ���jj�Zy饗��3Ϥ\��   ���  p�fgg��/:ɶ�Zv�   �d�p=s�dtZ���jO>|�p����.   �B�  ܷ������)��V�w��   ��;\�܍Vn�mV�_|��g�f���  �C�  �}9u���at���<6ҟB�    �K�P�c�9;6���ji�Zy뭷�cǎ���  ���  ��Ν;y��7�b�Z���k   ��J�B�Л�F'2�hVK��̡C����O  ���  ��g?���!t���R��y0���   ��)ybc;r���9��X=����#*��ַ  �� �{Ҿ>���ہNP�)������Y    ��J�8���̌ȝUt�̙�ݻ7���  �m�  �t�ƍ���ہN�>�������    ܻZ���7�sfl2�f+�Z:�g�y&   ���  ��~��ٴ���k/������   `A�zJٷ���c�Ѹ�Z�����������  �	� ����ѣ�����b��'6���    n�R�ޡz>�5�VK�������{��lݺ5   ���  ���]��s��:�c�2\�	    �7R��L��������_γ�>�bэ�  ��  �U�����-8�vo�͖�j    X:��*�;�̕���j�����E����n   ~C�  �V�����&V�C�l�   ���s���f+קf��O>ɥK��}��   �	� ���}�p��j��[����    �|��2;�ʭ�F`5���y��gS.�X   �;  �4�ͼ��K��6T-��
   `�<����c������F��W^y%����   p  ���fff&����R��<���   `E���<ގ�G'sw�Xi��y>����ٳ'  ��&p  �Ӆr�ҥ�j���9�e`�P   ��S-�#r�L��
��'Ndǎ�T*  �/�;  0ovv6G�	��R���mH�\
    +�����6����T�-�;+��h��_�?��?  X��  ���~>r��R($OlHū*   �j���g��oNV���hΝ;�}��  X�T  ��a�իW�����P�	    �oS�'�s�|6~7��Z�VN�<�;v���7  ��#p �unzz:���Z`5�����    �9��W3;���ə�Jj6�y�����0  ��#p �u��K����v���`=    t�]C��4�����u��ͼ��9p�@  ��E�  ��ٳg3::X-j=ytc    �\���щL��VҩS��gϞ���  X?�  �N����7���ޞR�o�O!    t�b!y|co޽>���f`�4��>|8?��  �w  X�<�Fõ¬��b!OnH�X    ��R,���9=:��V+�Rnܸ�s��e߾}  ��;  �C}�Q�^�X�B�����{J   �{���g��nLVJ���ɓ'�k׮T*�   k��  ֙���ǎ����2T�:
   ЍFj=�1��g�w+��]��������   k��   ֙�fvv6�vֳ��    ����j��\�򝑕s�ڵ\�pa~�  X��  ��\�t)�/_����Jv�   ��g���F3wf�+���_ώ;R.�]  `-�?  ���µ�jVZ���#�   `m(�}�yot"w�|sde4�9r$�7  `�� �:��K/��ݻ��V)��恔ڧ�    ���>�7���щ�5E�-���J�o�  `m� �:p�ڵ|��'���n��q{�T    kO�\�c������cǎ��g�M��#  �Ew  X��f:�V˂+ﱑ�T�z   �e��r���Ӂ�0333���_�e  ��Ge   k\�#���$V�#C�l�   �����J��|19X	/^̾}��u��   k��  ְ���|�ᇁ�����G�z   ���k����\n��V�+���g�y&�b1  ��!p �5�^H�����J)���   ���PH�m��{��j�.��{�nN�<�o��  ��;  �Qo��F���+�Z*�k�Sj�f   ����Pϻ��i���>Ⱦ}�2<<  `m� ���O�>XI�B!OlH��:`   ���^.���z>�9�VK���j�����K��  `m� ����ϧ�t0+kT�f   �l���P_%���,����������/  @�S  �s�ԩܼy3�����j    �7��W2٘��t#��ڷ��۷/}}}  ���  ֐������[��4X-g�po    ��3T�Tc�Ǎ�,�V���_~9?��  t7�;  �!/��b���+�R*f����    ��V*��p=��&�h���ƍ��㏳gϞ   �K�  k��˗���VJ;j����TK�    ��R/��?�9=��˥��u�ĉ�ڵ+Ţ�  Э�  �F���+�XQ{7�e��   �?lC����*�t�n`95�?~<O=�T  ��D  �5��^���d`�<8P˶�    �W��+�l�el�XN/^�O<����   �G�  ]nbb"gϞ���j9{6�    �מ�Z��_=��ri�v�ꫯ�駟  �}�  ��<�f�a+�R*�̓)
   ��U*��p=��&�h��e||<gΜ�_r  ���  ��G}�����JhG�_�<�j�    X�z��݃�|xkz~i��/���ݻ7�J%  @�� @�j��;v�+fT�F   �xk�<����;3�����~�ȑ����m  ��L  �.��+�dvv6��e�@-    �T��U21;��w���ʕ+�϶m�  t�;  t�7n����0T��ލ�   ��T(�w���F'3=�,��G���g�  ��  Ѕ^xᅴZ��r���yb�@
�    ��+ylC=�G'3�'�dzz:o��f���o  �|w  �2��Nn߾Xn��}#��;    ,��r1;����t`��={6���O___  ��&p �.2;;;�2+ᑡz6�+   �嶹ޓ�ٹ\��,�������J����  �lw  �"����\`�m�U��Po    `���eb����(�ctt4/^�Ν;  t.�;  t�+W����ˁ�V)����    �J*�G��ywt"s�V`9����y��S,  t&�;  t��^z)��
_=�7�G�    ��j�Bv���ͩ�r���������SO  �Lw  ��E��):,�]�2\�	    ���Z9��=�bj6�.\��dxx8  @�� @�k��gΜ	,������    V�ΡZ�4����,�#G��G?�Q  ��#p ���K/��l�S�\��    ������p=�Nd��
,�۷o��?Ξ={  t�;  t��W��ʕ+��T($�7��X    t�j��=C��c2��Z�VN�<�]�v�X,  �w  �`/��r`���П���C    :�p��m}�\��	,����������v  �Ρ`  �u���ܹs'��6�V��@-    Щ����\�g�K�>ȁ���  �3� �5����XN�r1�F    ���ճw��wG'�h�K��j��ѣ�����   �A�  �W^���l`���Sj�    �Z*���ZΎM�ڵk�r���<��  V��  :���xΟ?XN{7����   ��1T)硾J.O��R{��رc��O~  `��  �ü����a�l�f[-    �m�Ts{f.�s��499�w�}7  ���  �A.\������ri_���H    ��z�P�;�'�h
ai������\��  �j�9  t����\
�B�4�r�    �V�b!�����t`)5�?~<���w  ��;  t�7�x#��dX>��3\�	    t��ZOn�����l`)}�駹u�V���  ��;  t�����9s&�\�j=yd�7    �V�����\���Ri�Z9r�H~��  Xw  � /��b���ˡ\,f���    �ZR,${��9=6�f�X*�����g���  V��  Vٵk�����ˣ�R-    kM_O1��+�t�n`��W�O�8��;w�X�m  V��  V��Ç�?��r��_˖�j    `���ۓ[w�5�L����l�z��ɟ�I  ��%p �U��{�e||<��=����    X�
�B�������6���tΝ;����V��  �J� �*i6�y��7ˡPH�����    ָ�b!{�jy��T`����9r$�w  `�� `�=zt��SX���2P��   ��1\-�ޞ\��ݕ�s���\�~=�6m
  �2�  �
�����G���z%��   ����Zn��e��,��Ǐ�G?�Q  ��!p �U���/�_m
K��T̾��    �zT��yt���F'3�j���۷s����ܹ3  ��� �
�y�f._�X�R*    ֫z���*�p�n`)�Z��<yR�  +D�  +쥗^
,�����+   ��nko%�f�26�,�������{��׾  `y	� `]�t)ccc����Sʮ��     �a�`-�3�m�K�ԩSy�'R,�E  ���  V�ѣGK��ճo�?�B!    �(�5X�7�Kann.���/�g�g  ���  V�ٳgs�Ν�R{x�7�՞     ���Z9��z�O7Kᣏ>�7���j�   �C�  +��lί��R믔��`=    �o�s���ىܝk������^�_��_  Xw  X'N����L`)�<>�?�    ����Bv�r��T`)\�t)7o����p  ��'p �e��Ϟ=Xj��{�W�Z    �P����=�br6��?����  ��  �ّ#G277XJ��r��    ܛ���uw.�s��b�����իy��  ,-�;  ,�;w��O>	,�R���7    �w�B!{�j9=6X
�����  ���  ���Ç�j�Ki�p_��b    ��3P)塾J.O�kbb"~�a}��   KG�  ��ڵk��/KiC�'�j    f{57g��m��7�̞={R,% ��"p �er�ȑ�R*�ٷi     ��
�ޡz��H��,���lN�:�o~�  ���  ���r�֭�Rڻ�/Ւ     X�z�8�������b�>}:H�,� ���?k  XǏO�e��������}�     Kc[oOn�m���\`1��f^��<��S  O�  K������T`����ytc_    ��S(�g��S�'ҴW�"]�x1������   �#p �%�^ii����R*    XZ�R1��r��t`1ڷ����k����  `q�  ���|������ʖ�jF�     �ckoOF�gs{f.�W�\���x  ,��  �H{��̙3���S*fφ�     �k�P=�\�H��
,T{���������   'p �%���[ogI��ЗJ�    `y�J�l����Ÿv�Zn޼����   #p �%�h4r�ܹ�R�W���    `el�dt���ٹ�b�Wܿ���  X�;  ,�cǎenΡK�T,�ё�     +��ճg��wG'�jlttt�	  p��  �H333���Keφ�TK�     +��\̃��\��	,F{���?�a  ��'p �E:r�H��f`)�z���    `ul�f�n#S�}Y��7o�/��֭[  ��;  ,���T>����R(
ylc    ��S���3T�{����x�����O  �?w  X�W_}�z;Kf�po�=�     �����m}�\��	,���x.]���۷  �ww  X�;w�����0P-g�`=    @g��_ɍ�F�猜�p'N�� �}� ����+��Y�B!�F    t�R��]C՜�
,���d>����ٳ'  ��� �ܾ};��y
�B`�����    ��U���ۓk������/)p �� p �x��K��RΎ�z    ���p57��ef΍�,���tΝ;�}��  ���  p��_��/��"�X� �؟��     �c������܍��B����w  �Gw  �O���j`)<4P�`�k    t��rFj=��,���LΞ=����  ���  p�����Ū���9�    �;����L#�f+��N��_q/�  ~7�;  ܇#G���rx��=:ҟR�    �;���_���w1;;�w�}7�G  �w� �=���Os����bm�W2��    t����\�j���\`!Μ9�Xq ��C�  ����_,V{�}�H    ��S(�k��wG'�h4�� � p �{����֭[���9ܛj�2    t���b�������B�>}ڊ;  �w  ����Z`��zJyh�    ��=�_͍�Ff����������  ���  �\�v-7n�,֣#�)    t�R���k���T`!�  �	� �8v�XZ-+<,ζ�Z��=    ֆM�r���rkf.p�fggs����߿?  ��$p ������,FO��]C�    ֖]C��s�N�6RX�w�yG�  ���  ~��G�Zog�vo�OO�    `m��
y���Kw�����LΝ;�}��  �/w  �n޼�/��2�C��<�_    �6=�_���l����j��� �� ���ꫯ�������     kW�;�#ռc*p��������G  ��  �[����/�,Ǝ�����    �m��rFj�N7��ԩSw  �o�  �[���[�V`�j�b�    Xv�rkf"��o�ܟ����?>�w�   p ��cbb"��y`1�n�O�X    �>���_���Ӂ����o� ���  �9r�z;�2R��?    ���@oO������\�~��w>���ر#  ��	� �i_z����B����    `}�9P�����:y��  "p ����W_��΢l��^.    X�*�l��s}����+W�d۶m ��L�  �6===�',T�T�Ã�     ���Ռ�m�iO��t�ĉ�˿�K  `=� ��;v,�f3�P�7��T,    X��c�U�ٝ����իW��  �+�;  |eff&/^,�`���}�     �=�_͗S���3�����/~���� ��J�  _9~���v�P(d���     �F��Ǉk���T�~ܾ};_~�e6o�  X��  �{�����z������+    ��X-g�����F�^�Z������ ��H� ��w�ĉ����T,d�Po     ~�G��5�H��g7n����x  �� �u�ܹs��j��R1     �M�\��z%W'g����������  Xo�  �k��^ff*�0�=�<4P    �ﳽ���ӳi4͸s�^�:�Q�T  �� �u���,Ԟ})    �{�����������j����������  �z"p `ݺp�B&''1R�dc�j    po��˹6U��l3p��g�g�b�  X/�  �['O�,D�PȞ�}    �W�B!;k9=jx�{�l6��;����F  `�� �.]�~=7o�,���z��R     ��@O)#�rF��{u��Y�;  �� �u���ぅ�)��`=     ��@57�6�l�I��ȇ~�G}4  �� Xw&''s�ڵ�B��؟R�    �����y���Kw���;�#p `�� ��=z4��i�_��-��     ,ƃ}�|19�Y3�ܣ�x��˗��C  �:�;  ����l>���B��M�`�    X��%�;�9k:p��z�-�;  �� �u�7������Sg~��_��g8
IX>���wk�)W���S�����ڿ|�U�hW�lY�@� 3�l�ȑ% �������K��t�G�;��n�i]��.    ��p�V���vl�{f�ɼx�"���brr2  `�	� ȍ,l���	8�l�=[o    8K��VㇵV�I]�~=����=  `�	� ȍ�7o���^�i]��c���	    8[�B������ĳg�bgg'��j  ��Rh  ��}�]�i�Iį&    p>��w��������;�����o�  0��  �������	��ǣ���     8�R!.U
�|g?�$?~�n7�Գk  ��� �\�������*��d�     ���F+���6�9�l���o��/��2  `	� z������pZ��ע�&    p�*�4>���ik/�$��k����ي;  CI� ���ӟ�pZ�b!��T    �"|4R�������q�x���q�������  ��� �����+++����z���v    �bd�I~8R�ٍ����s�� ��$p `����G�z�n8��J)��+    p��k�Xj����g{{;���bzz:  `�� Z�n7fggN���     �h٩��Vbf};�8��ύ7��c  �0� 0�n޼�N'�4.��1^-    ��p�Z���B4�<��x+++�����SI w  �֝;wN#������    �ٯF+q{�pׯ_����:  `X� JO�<�V��N��h-�%�I    ��5Z.�d�k���y��qt��H�4  `(7  J��N#M">�    @?�d���N�z����t:q�������  ��� ���-������G��(��     ��^�V���cŝ�ݾ}[� ��� 0t���?Y��T
i�Yo    ��ߍVbmg?<��8;;;������  �N� �P�v���ѣ����z;    Ї��4.�J����6��ύ7��c  ��� 0Tn޼�N'ऊi�V    �}<R��;��ur)�XYY���ݨT*  �L� �P�s�N�i|2V���v    �OU
i\�c�eŝ�]�~=����  �A&p `h,,,D��
8�,l�h�     �죑J,o[q�x�?�n�ij� ��%p `h���g�i|:^�B�    @?+�IL�K��x�N�w�ލ�?�<  `P	� 
�r���J�Ie��^�    � ��Q�g���Xq��o�� 0��  �?��O��P�S�t���v    `@�$>h��ɖw�ngg'���bzz:  `	� x�n7=zpR�z�t�z;    0X>l�c���]�/-�q�F��  Dw  �_����t:'��Ɇ�v    `��$�5�1���6+++������  �� ��w��퀓��
q�z;    0���˱�lǞw�q������  �� ������V+���D#     U�D|8R�ٍ���y��q  � � 0в��^�J'3Z.��z9     �t�t�������������>  $w  ���~,--�ԯ&�    0�V��x���6�o�� 0p�  �o��6�]�4�L��~�f�    Wk�Xh�Yq�^�x�f3�F  ��� 0��ݻpR�Zo    �H�D\k��w�q�ƍ��o  �� ��������'�(b�z;    0dVܷ�����277  0H�  ��ׯG��='�	G�    �'�V�G*1��p�N���ߏ�>�,  `� 8�v;���N�^*�T�     �h�V����س��[ܾ}[� ��� 0p����;��n�I��x-�$	    �a����(���n�Q^�x�f3'� ���  �{���D�X���J     �j�x�lǾw��ƍ��7�  �;�;  eqq1���N�Ӊz�n    �]!M�z)��G���  w  ���ף׳@���4���    ������9B�Ӊ����g�}  ���  �v�KKK'�w��H��    @>�w��Iӊ;G�}��� ��'p ``ܸq#��n�q*�4��     ȓ�x�jG׈;Gx��E4��h4  �J� �����	8�O�k��   ��)�IL�J�p�lP�o�	  �Ww  ���b�Z���d/p��T     �>����~t{f�9���\  @?� 0�_�p��׭�    ����\��b��8L�Ӊ����g�}  Џ�  ��v�KKK��^�|h�    ȹk�R,��aÝ�ܾ}[� @�� ��nܸ�n7�8�ף�Zo    �RH�J��Z{���؈f��F#  ��� �{333�)�I|d�    ��G�J,����s�^�w00��7�  ��;  }�ٳg���p�Gk��    �W���T�+�V�9ܓ'O  ��� ���������$I�[o    xՇ����#������\|��'  �D� @��v����p��F%*�4     �?�b��b�h�����w  ��� ��u����t:��d�     ��Ñr�X�s�������45" @�� з��8ΥZ)�B     ��r!�B4���^�w�܉/��"  �_� �K�v;�����w���    ��Z�3�������  ��;  }��o�=X��-c�R
     �6U)�\!�ݎ��l\�F#  �� �K���8�'�     ��$�F%f7v��%��_�5  �� �;ϟ?�V��6�b!��+    ��֊1��D������w  ��� �����瓱j     p2�$��z)�������ӧO�ڵk  �� ����ɓ��)�IL7�     �q�Q��V;�F�9ĭ[��  ��;  }eff�`%�棱Z�$     8�l<�r��Z�������v���i  ��$p ��d� �6�1��Xo    x���X�ޏ^ό;?���w�ލ�?�<  �}� �7��v������H%J�1     �VLc�\������	� �w  ��_���1���Z     ��>l��jss3Z�V���  ��E� @߸w�^��\iT�V*     �n�\���][�N����׿�W_}  �� �kkk����6��    �Ƶz9^���c�;  �� �������h�c�0     g�R��B��n��vwwcii)���  �u  }a~~>�m>�     g#I"��J1���[�n	� xo�  �w>�v�p�R!�+�;    �Y����Is7����y��Yt��H�4  �	� x����p�i     ��b�ĥj)V��^��t�>��  ��&p ���?�8JvL���     ��Z�,p�Pw��� �^� x�~��ǃ8ʕz%*G�    ��F1��r!6۞��s���CEi�=  K� �{������G��     ��L�Jw������~���  \$�;  �M�����p��r1�*n[     ��T�s[���t^u��=�;  N) �{s�Ν��8�G��     �|%I��Z���j}}=����X� pq|� ����R*�q�!p    ���R<i�F�.����|��  E� �{��}����Ñj�I     p�i���X��x�����  \(�;  ��_�������p��k�6j�    �"]k��ass3��v���  �� p མ��	8��z%*�4     �8�b��Bl�;/e�E�oߎ��
  �w  .\����ŋ��|4f�    �}�����ѣGw  .�� �w��̓�8�H��R     p�j���j�n��R�ٌ����V�  p��  \���Z     �~$���K1���R6\t�֭���/  Λ� ��j�bcc#�0�4���r     ��\��b~k7�ʫfgg�  \�;  ��͛G�n���$    ��SJ��,cuw?ढ़����܌���  ��$p �B=|�0�(�Fk    �����yU�׋۷o�W_}  p��  \�lգ�jf�Z�F�     ���BTi�t�/���	� 8ww  .̍7�=�0�F�    @��R+��V;ढ़��X__����  ��"p ��<~�8�0�4���r     �?���1�l��^u�֭��o  ΋� ����������Q�B�     ���&1Y.���~�K  �I� ���y�f�Q��V    ��3�(�������a����  �� p �B<y�$�0�R�K�     ����Q-����dz�^ܾ};����  �� p ��mmmE��
8̵��     ��J�s[퀗�>}  p^�  �����/�)�iL��    @��Z/�|��^�����������  ��&p ������F%
I     ��R��d����/ݹs'��_�%  �	� 8WقG��8̵�j     ���e�;?3??/p �\� 8W�n݊�3K9�D��R!     ���BTi�t��V�u0tT�� �l	� 8W>8̵�    ɕZ1���l��~�?��  gI� ����ߏ����ו�$.�+    ��Z/�|�n�G�	� 8sw  �͝;w��uT)o�nT#M    ����L���������<<*%H  ��. 87���8���v    �At�^��3?��c����}  �Y� p.�������׍��     �g�R<Xr���2<� p�T%  ��l�=���u�T    �����\+��f; ���~�N(M�  �� p �\d�Q��W�     `p]��^�w������&  �,� 8Ϟ=x�T�|pt-     ��^L�־�\�333w  Ό� �37;;�N'�u�#�     `�e+�����  ��"p ��ݹs'�u�4�K�R     0�.�J�xk7z���᣹����O  ~)�;  gnqq1�uӍj�I     �R��D�k����w�
� 8w  ����R����n�Q	     �ǕZI��O�={  p�  ��[�n��^*�h��    �0����&���t:��!����  �_Ba ��ZXXx�#�     `��IS�b,m;ٕ���?� ���  ��f�;;;�J�$�6*    ��R+	��ɳg�  ~)�;  g��x�D��B     ��r!��4Z�݀l��jE�^  xWw  ���Ǐ^��H5     ^�k�x����w�^��?�c  ��� p&��n������&q�^     ����We�Hw  ~	�;  g������^u�^�4I    ��UN���c}w?�ŋ�Hi�  ��;  g";n^7=R	     �_��.p'�"���ŧ�~  �.�  ������WU�i�WJ    ��"M"�{�o�߿/p ��	� �����boo/�UW���    �$1Y)��+�D,//  �+�;  ���۷���W]i�    ��r�$p�@�ݎ���  8-�;  ����|���B���n     ��x��4���Q"~�����/  NKq �/��v8�UW��    �N�$1Y)���^��'O�  ��;  ��ݻw�׳���	�    ��r�$p������PR��  �!p ����	x�h��b!     ȟ�r!Ji{]�8y�$=z�(~��_  ��� �_dyy9�UW���    ��R�K-+�Dܿ_� ��	� xg+++�����;    @�MUKw<�<  ��  ����.�U�RT
i     �_c������N7ȷ���X[[����  ��� ��^u�z;     s�R��-�;w�ލ���*  ��  ��v��f3�$I�J�     p�V���� �I  ��� �w����G��xi�R�r!     h�
Q-$���.!�Z�V���G�(S �d|s ��<x� �UW�     �����x�l��&�������  ��� �NVWW^J����;     ��r�(p����� �� pjϟ?�N��ҥj9Ji     �R�X�z��=��nmm-  ��  �������    8�TE�N���^lmm���H  �q�  ����B�Ki��T�     �Z9��333�?�!  �8w  N������F�K�b�$     �u�B�b��n�oO�<� p"w  Ne~~� r����+     G���e�=�^�x  pw  N�޽{�ʎ�    ��\���=�:�N<�<���  �F� ��,--�4^-E��     �Q*D���n�	�y�)	� 8�� ��v��l6^�R�     �R�O�V��nqq1  �8w  N,[���z/M��     Ǚ�܉���:TJS�� p4�;  '������F+Ũ=�    �x��4Ji{]C:y�)-,,��  p�;  '�����e��     �P�$q�Z��������  ��� ����9����J     �IMV
��
rnyy9  �m�  ��ݻw���L��F�T     8��r1
I�r��j���~��%  �"  '2;;�ҕF5     �4�$b�R��;�A�=|�0~���  F� ������4U+     ��T�$p�`XI� �Q�  kcc#���2�Bc�;     �7Q)F�Dt{A�=�<  �(w  �����G��I3��r�     �.��}�\��]+�y�+���D�Z  x�� �c����t�^	     xW��{�e�J333��_  �N� ��^�x�)�i�WJ     �j�Z�d#�ٱ��,	� 8�� ��Z\\�N�����"I     �Y)Mb�\����y���  p�;  o�	/M�+     ��d�(pϹl`��lF��  x�� ����!��g��    �/5Q)��f�c�^/�߿���  �*u
  o���������     �T�X�j!��N7ȯ���;  o� p��������L��     ge�R����=ϲwQ  �:�;  G�w�^�Kw     ��d�K�� ������nG��  �G� ���<y��Ҩ�
     ge�\�B�D�����Ç���.  �%�;  GZ[[�L�+     g)M�-b}w?ȯ��9�;  ?#p �P�V��XH�\��     ��d�(p�9�K  �N� ���ݻ�I�����    ��7^.�����n7�4  �� 8���|@f�Z�B�     ��j1�Z���� �z�^<~�8~��_  d�  �����K�r     �y�(������� ��;  o��ۋ����̥Z)     ༌��x����J  �Kw  �p����L�T88     ��d��ͽ����|��ގn�i�  � xCv$d�j�     ��$��������bqq1>���   �;  oX^^�L�J     �m���	r�ѣGw  � ������H($I�W�     ���#��_nF�P��   /	� ����كc ![oO��    p�j�R$흿������V  @F� ��<|�0 s�V     �(#�$��^$�Wr);e����155  �� ��YZZ
�LV�     \��F�Zތ��� �<x p @� ��5�̀Z��b     pQ��5��pA��c��  �� �������0Q+     \�4Ib�T���ݨT*A�lnn  � �Iv�#d&+w     .��1��E\�z5ȟ�����ىj�  �� ��<{�, I���
�    �xY�~s�iLMME�P�gvv6~���  �%p �'/^�)�TH     .�d��b!677cbb"ȟ���; @�	� 8�����`�    ��%;etz|$��������Z  �ow  <z�( #p    �}�6>�W�c{{;j�Z�/��;  �&p ����\@�$1^�    ��d��{u�݃����   ��  X^^���&     ��h�#�r4���t:Q(�|���� �� �[[[U��     �L�������܌��� _�={  �� ��P`R�    @�9�766�9���  �� �x��a�z� �
I��;     �_�����ۋ����jA~���F�ۍ4M ��� �����R$     �_�T��F-֚�+���y��i|��G @�� ���Հ���v     �����A��l6���D�P�cnnN� �Sw  ��jL
�    �#�&F㇅���z���A~���  �$p ȹgϞE���RH�^r{     @��:6i�D�׋���{�lmm  ��` ȹ��ـ	��     ��b!���z,o4coo/����V��������(�� @�� rnqq1`�"p    ��d+�Y���V����5����  �E� �skkk�    �GW�?���lF�ӉB�����  ��  9��vcww7ȷb�D��     ��+��H�$z������A>���  �#p ȱ�X��a0�6^)�     �~S.b�^�������i�Z @�� rl~~>`�Z
     �WW�?�{{{����j5~�i��j���h  �w �{��Y�X�m     ���X#~|����Y�,pϏ�D�/��"  �% @�e�ɷB��H�m     ������~��ڊ˗/G�$��3� �?J ��ʎt̎�$�F+�H�      ���ʥ�Vbsg����G�ٌ���`����  �"p ȩ'O�D���m�Z
     �wW�?��Z�{>���  �"p ȩ,p���[     ��ձF<x���ϭV+:�N
�`�e��Y�^�V �|P�  ����r�o�߮��w     �ߕ�7�ڳ����`�e'����o~�   �  9�����h��4	     �wc�J�ʥ�n�����=?�  9"p ȩ��N�m��v     ��qe������s�ݎ��ݨT*�p[[[  �C� �C����9�o�R     ���2���=���܇_��  �C� �Csssc�;     �cz|�ϲ�}jj*�$	����^t��H�4  ~w �Z\\�^*D)��    ��1Q�F�X��~�ϲ��jE������R\�v-  ~w �Z__�m�j�    �����_m�����>�V���o~~^� �w �j6�A����
     0x.���ܳ��N'
�B0�VWW �|P�  ������C^�m�b�    ���-�fkk+��ǃᵱ�  ��  gfgg����UL���     �A35R?����M������  �A� �3O�>�m�\�$I     M�X��Z%6�;g�s�ݎr��l�i}}=&&& ��&p ș�ϟ�6Z)     �K#�7�L��>55���y�; @� rfkk+ȷ���      ���z<Z^{�����}�-//  �O� �#�n��xN�m��6     ��55R?�������ىj��/^  �O� �#O�<�^��W��F��     �K#�H�$�����V��ë�j  �O� �#Y�N��VJ     �,��'�x��f��/_�S�ӱ� �w �YYY	�m��     ��wy�~h������Q�Ղᴰ����� ��n ȑ��� ��*n     |S������d+��ᵼ�,p r� �Ɏl$�FJn     |S#�#��/_�$I�ᳶ�  7u @N�������k�\�B�a>     �o�V�r������v��j���h�'�  7�; @N<}�4ȷъ��     �l����桿�"h��p���  ���  '�|-��    ��x[��l6���E�8�t�d�����r9  N
 ��X]]�m�R
     S��#���Y�>22������O ��$p ����moIz���|�dI����K���Z ȓY�=c�߻�lk3�̮mI�DuU� �)e��BT������A��� �:      ?\�}������� �M� P��b��b2��    ���hg�qܯ7_����H۶QUU��_�5  ȗ� � ���v��u>��    ���?�}3p���qA^�u~  �r (�O?���|�?     ��>��~���w!��=?��2  ȗ� � w�Fu     @n���{�E4Mu�<'���ݫ��   ?w �|��1(W5�\�    @���揾���>޽{�c��?<�ۿ�[  ��; @>����ۻ�     rs6�d4��v������	�3���?� 2%p (�r��uf�    ��]�g��͗o�{���mۨ�*ȇ� �%p �\w`�^��r�O|�     _Wg������������˗   OJ ��Y��|�k?     �z6{�=���V�   OJ �����wP��Q     ���'��"��}� ����&㪪 ��� 2g��l���Q�`    �|]ΦQ����|O�w����Y��O�>ŏ?�  �E� ��ϟ?庘�     rVU���O����w�w/p��_��W�; @��  ��k)���     ����ٓ�n�}0y�� ȏ�  s��:(��H�    @���G�Ӷm�V���/i���	  �#p ������	庘�     r���i�z��D����  ȏ�  c��_�r�*&u     ����E������?y�n� @~�  ���cP��q     P�Q]��tw��w��4����t:���d���b8�@ �ķ; ��}��9(����}     �q=�=�w�w�{�������  �x �ؗ/_�r	�    (���,��G���>|� p ȏ�  c��"(�|X     ��j>{����ml6���A�nn��  �"p �Xw8K��#�;     �x7�<��݊��=n4 ȏ�  S���~��4�QW�     �R\L'QU�h�ǟ�t����u�>7 �G� ���~�I�^�ٰ
     (I��O�q�\?���z��.�C�L��h ��� 2���?�:��    @y.��'�n����2H[�4ѶmT�� �\�^  2�믿��     �Ҽ�M��?o����b!p�D�\�Ç @�  �����5�    (��|���.�����1��}��Q� ��; @����5��    @y�=#p���.r���A�~��   � �L���L�j��    �Ҽ�Mٻx�)����p�1 @^�  j�6��	�t6�5    �2�*�&��[m��~7���� �� @�>~���e�3�     �z7�>9p��v��lb<�r�1 @^�  ��矃r�-�    P���4�߯�O~��-pO[��
  �C� ��_~�%(�|T     ��r6y�������*HWw����]���  �� d����A��F��    P�w��޿\.�mۨ*2)�n8� �A� ������Lê�q�     �r]�=/p�t+���}��)��?�#  H��  C��*(�|$n    �l����x����?#pO���M  ��; @��ۧؒ�����     p9�>;p'm>C �|�_  2ӭ�����L�Q     P���$~�����o�&��uL&� M�� @�  ����SP���     �b6}��t��tm6�   w �����A�f�*     �t�����>����4u+�  �A� ������\ӡw     ��=�}�^?D�u�=U�
�|>  �&p ����]P�I]E5     ��l2��`���Y?��A�����  �� dF�^��Ȣ     t�A��x��ͳ~n�\
��������  �M� ���j�i6�    �o.��g�݂;麽�  �'p ��f�Z�1V     ���lq�i���Y�x<��c �<� 2���2M-�    ��:��/�K�{�,� �A� ���j��>(�l$p    ��\L'�\I_^^�q�1 @�  ��_�r�,�    ��:��w�ݠ�`0Ҳ�n ��	� 2"p/װ���r�     ������.n_��1�N��4M  �O� ��ϟ?e���      ��hX��o�����s��.pO�b���|  �K� ������L�Z�     ��|6���ų��������t7� �&p �Hw�J�f�:     �?��N����z���m��̤�������� �t	� 2�]�I��#�;     �����������Z�,�'�˗/ @��  �l6A�,�    �?��M��nXH������   mw ��4M�if�     ������}�Xć����  }w �Lt�d�m��b\     ��������n��ƅ���LJ��u  �6�; @&>~��i:�b0�    �?��GQWU4�uk����A:��m  �6�; @&>��iRW     |��d���V���q�1 @��  �����4
�    �[f����b�e���f���x  �I� ������L��     ����C��n��6F�Q�������� �4	� 2�Z��2Yp    �o����ӗ˥�=1���w ��	� 2��R��Ђ;     |���nd�ݻwA:�E  �.�; @&6�MP�qm�     �e>9~������  �� db��e��    �������n��e6��� �6߼ 2��R�z0�a5     ���&��j����� �� @��  �h�6(�dX     �m�aú�]s����r)pO�z�  �%p �@w�����L�U      �7��vyx�l<-n> H��  777A�Ƶ�     s6�o6�h�&��ͪ)� �M� ����۠L�;     <j6�;��u�����?F   ]w ����e�    ������r)pO�~���m��<G H��  �rM�f    �1g��ѿc�Z鸿�����   =w �,��L�a     �����/����e��`�����  Qw �X)פ��     �����{�w�df�Y�_�|	  �$p Ȁ��L�`ue%     s69~��#pO���]  �&�; @v�]P���z;     <Ũ�^ۦ9��,�˸���o�X  i� d`����w     x��x��q��[u�� H��  m���    ��M�]&�>�w���X��1�L�~�>'  �$p H\���4�     <�t�2��r��'��  �� $���&(Ӹ�     x���e2��j��v�  �$p H���]P&�     �t/��^���s2 @��  �[,A���*     ����F/�{v���k8�����  ]�i $�5���     O�R�n�]��o��>  H�o�  ���k\�     <�K��󙳳���,� ��78 ��	��e�     ���鿻�����
  �"p H��2ՃA�w     x��^p�����  Aw ��	��4���     ���0�jm�?�w����l61����  i� $�;<�<�     �y&�a,7��]����ߺw  �#p H�v�2���eTYp    �皎^.p���/..���� �&�; @⚦	�3V     <O���t�u+�  �G� ���n�gT	�    �&/�o6�h�6*g���}F  �G� ������k��     �\/������t���  Mw ��5M�gT     x���W����Ƕ�m  ��; @�,��iT�    �^:p_��A�v�   =w ���V�\�     �y&���N	� �$p H�b��T,�    �s��/; ��M�Dm����  i� $���>(Ө�    �s�^!D�V���΂�i�6  H��  a��2(�`0�Z�     �6�|*�^��=��� ��� �X,����     p�q]����w�ɂ; @��  	��^�Z�     뇛R_r�[��o��&��q  ��; @�V�UP�a���2     P�Q]�f׼��k���U�u�?�`��  -w ��u��gX�p    �C�������l6������  �!p H�n��c�     7z����z-p�)�Q  �� $L�^�ڀ;     �[pi]�N?m��   -w ���m�gd�     6~�w+��� H��  a��44�     �^'p���18���  �� $�i��<u�p     5z��N�O&��_F �G� ���m��*     �Ì�����k�{Yp H��  a'�Tp    ����;�#p H��  a��4��     {�w��` @z�  	��iX�p    �C�ւ�����  �� $L�^&�     p��+-�����n�1���h�&  H��  a�A)��     ��R���V���"p H��  a�2��    �p�+ޔ��l�~� �G� �0�{y�AT�;     jT�^��-��/w ���  !��    �8��Ҷm  ��; @���8���     �y��}��=,��u��  =w �D��L��     �RW��6$��n�=���  i� $j�Z���     p�nPf�J��f���t�w ��� ��R�     p���b�J�g8�"p H��  QG�T�p    ���A�_�wo��   'p H���LU      Ǫ��;q��_��}  ��; @������     G{��}��E۶QUfk���,  H��  Q��(�w     8ְ~���*�L&  <��  Q�&�$p    ��_y]}���{b��
 @r�  ����Ay*g�     p���;��� @z�  �j�&(Ome     �&p ��� @B*�;     �~�+S��m   �� $ʂ{�*};     m���]���c`��ڶ��?s  ^��  Qݡ(��     ǫO�(�E��$x{w ��� %p/Sm�     �Vׯ;o6�{Ot�;  �� $�i��<�    �x��4�;�`8
  -w �D9�+��     �w�=��v��( ��� %p/���;     �7�Zp��; @Z�  �j�6(��     �w�A��� @Z�  ���^*�;     ��{��E��(x[�� �E� �(Ke:Ţ     �:�y���<W H��  Q�&�$o    ��2p��5M  �C� �(�;     @�	����; @Z�  �rW�S-�     @�':o��v��3 ��; @��     ��N�[pi �t� e�     ����� @Z�  ���^��DW�    @�N4��Vw��u]o�s5 ��� � �T>w     8����2݊���mYp H��  Q�2Yp    ��:p�N���� �E�       @QN9'��  ��	� UUU      �|Չ�y[u]  �� $�Wg���     �6��p @Z�  ��     �����y� ��; @�,M��,     �7�6Mm�z���  �!p       �Wԭ�O&�   'p H���2���      �Ӟ��]����C� @J|{ H���Lw     H�n�ގ�j  i� @BZ�;     �����&  ��� $��D�ڶ     �8��1Ղ�۪�:  H��  Q�2�-�    ��N}�.p[w ��� 5��w     8���� H��  Q��Դm      �i���m�>�<�y��  �"p H���2�-�    @����x��?,  H��  Q��tq��e      Go1(#p;áD
  %�� $���,Mӄ�     ��{2]��۰� ��; @�,���;�~�E     ��[-�  �� $��Dy��     p��8m���n4�s5 ��� � �<]��
�    �h��a<  =w �Duk���7     ��V�  �%p HT]�AY,�    @��  �4w �DUU��;�v�&     �-eڶ}xy�  �'p H�p�\i���     ���jP�������   -�( �D�F���A{��w     H�����  �� $j2��x���f׶     gۼ�y{�sZw ��� %p/�o�w     8^�
�KQUU  ��; @�\_Y��ܛf     �q��� ��; @�,���w�     p�]�6�2�ӳ� ��; @�������~oѻw     x9��Q�u  ��; @��M���}��    �X����v���x� ��;  $��;     ���}�r�'p H��  a�� ���9����	��     p����w�{]��i��  =w ��u�������     �X����� H��  a݂;e�-pߺ�     ��ց;�3ʣ  R� @ºw������b?     m��K!p H�op  	s�b~�ݴ�      ��{�A��n���i  �� $̂{��[p    �c�堌�Ӳ� ���  fq��?�~�+S     o9(#p?��h  �E� �0�{����,�    �Q���]�~Zw ��� &p/����     p��ݿ����I��( ��� �0�{������     R�Xp/�x<  �"p H���������òL]     x>�{YF�Q  ��; @�\�X�<�����+�=     bۼm���t�6��1�S� �G �0W*��������Wy     8�f�{��g���Nc:�  i�M  a��$��?�]w��    �C���{g��	�Od6�  i�M  a'��]Qڽ~��     �����i  �� $́\��v�����;     ��C2��QUU  ��; @�\������C��֡7     �C2_;���u�;  �� $���,�����V]     �`������Ӱ� �&�; @���σ�}u�}'p    �C�a��1fsu]  �� $l:�y�z����     ��m�����OC� �&�; @ºk��C�|}�][p    ���aHƳ���F @z�  �A����?�߶�-    ��m,�C� �&�; @��F𜭯po-�    ��6۷_p�l�4�  i� $n8�v�����}-p    ��m[��� @z�  ��w�e�     ^�~���9���4&�I  �5 @�\����povw     8Ķ�GX.p?�; @��  �����M�~�`     ��mv�苦i������f�   =w �č�� _�Zp�O��|�    ���4�YN��_�t:  ң� H��=o���;     <W�ܿ���3�� ��(b  7�L�|}�p{�k�<     ����l���uvv  �G� ���l��{��mf      �M�כ�	^�t:  �#p H��=_�������l     x��?���_�`0��� ��� 'p����[V�    ���tC���uu�;  i� $n>�y����҂;     <�J�^��  �� $�ݻwA����7�me�     �m%p/�p(� H�or  ���fW,~/�&M�;�^	�    ��V�b� �� @�+��	����m      ϳ���|�x��L& @��  �(���n����     ����c��g5]�����i  �&�; @F�Q��� /�_p�    �s���^E�m۟�>G��<  H��  ��8���ٛ���n㡯�     �}��[pUggg @��0  ��fA~;����     �4��� ҥ� ��t:�����r��w��     �dݳ��m���\\\  i� d`>��y�`�o�     �g��ryy  �I� �yz�`{��     �4�r��� @��  ��鱃��F�     Oշ����\9\UU @��  p�b�]p���      ��o7�Zp=w ��	� 2��ݻ ?��[�;     <U����g4  �� d�[��^�����{��f     ���x3j�l������ @��  �����}��    �S�q8Ɗ��L& @��  ��(v��-�p���`a��     ��vMۿ�\��:��i  �.�; @&�C_�r�ءvw���b2��    ��,��[o︝�u���   ]J �L�f������Ֆ��F�     ���魨�_���y  �.% @&&�I�����ϭ�     ��,6�\p���; @��  �p�b~�r���+U    �O�=�۶^���e  �.�; @&,Q�婋-��^�
     }�<�,ggg @��  �x��]P�;�     �����?u���QUU  �.�; @&�����,zz�*     ���r�r( ���F �����?,RX���S?�Ū��3     �ݙ�b����s��7� ��	� 2�]�ؽ��	���+U    �/V�]�B�b�f�   mw ��tW.
����w�ӑ��     �5�M?��;�_�|>  Ҧ� ��d2��z��9�݊��     �n��o���;??  Ҧ� �H�Hq{{��;���     ����+�/���2  H��  #)���w     ���%y��}  �6�; @F...��,�     �M���_���u  �6�; @Fؕ��     |���PL)�ATU  �M� �W.��9�-�    ������[pY��(  H��  #WWW�C�r�^     �Ϻg&��.(�x<  �'p �Hw�b�j�&H۳���h�6jWn    �tg�mk���$  H��  3�Ջ��t1�b����C[     ��/�~߂�Vޗuvv  �O� ��n�b�Ze���     �G��MP����   }w ����󸹹	���Ŗ/�u�u      �c��,��� @��  �q�b��~@     o��yY��� ��	� 2��ݻ }-�     p��D�YpY�׮� ȁ�  3�)�0��~4     ������y9UU=�  H��  3>|�sg�     �`���v�D�=w��o��:  ȃ�  3�������,ˮmc���l<
      ��O�/g<  y� d����ߋ$|�!��A��     ��n�	�1�� �<� 24�Lb�Xe�[��O��     Hc���sqq  �A� ��n�B�����-�     �oR87?�y _wuu  �A� ��n��ӧOAY,�     ���n>�?��c  ��; @�����/�KP���*     ���[[p/ɇ �<� 2��?i;�@ۂ;     �ݮmc��e��*�C @.|� �п�˿�Yow��51�     %�[�1
c��e���   w ������~����n����<     �dw�MP��t  �C� ��n�b�Nc���#p    ��<��݂��8??  �!p ��l6��v�
     (���yyI��� �|� 2uvv�?�t�b���5     ��}������Ç   w �LuK��_�����2     �t����?  �� d�A^�n����_     (�r����	��=��� @>�  ��ӟ����@}׶q����t     P���:Ra��x��(  ȋ�  S�����ݚ7e�Y,�     �f�
�1{& ��; @Ɔ�al�� =�,�t�~     P��e:���㝟� ��ٻ���3��/ �)J")q�,K�▇�޻�\��]՗�T�S��$�'�<E�e��'� �igQ'qEX�y��w�<�������� ������sh�2     9��W������d  �_�  }l||<vww�lJ���v�����j     @^m[pϕ�g�  �E� �ǒŊ�ϟ�����w     ��lF� ;��
܏off&  �/w �>f�"ۊ�b�Z�#���f��clh0      O�*��I��x��'  ��� ������u�Ֆ��}�;     ��]�V�n��xJ���H  �	� ���=ێs���ۏS     y��d���x��� ��#p �c�bE�\�l6��9�Q{�R     ț�j-����񌏏  �G� ��FGG�\.�s��=cO�    �Iض��+gΜ	  ��� ��MNN
�3�8G�-�     �L�Պ��zd������� ��#p �sgϞ��O��s�gI�덨5�1<P
     ȃ�j-��vd�q������  ��� ����l�M�]nٮTc���     �<��ۏ,��~<� 066  ��; @�[XX�鸇�M�;     9��ųD�~<CCC @� �����(�J�l6�l9��     �"kw�d��w7>>  �'�; @���D�R	�币�Fe/      /6-�����T  П�  9p��)�{w�e�\�V�Er     �\����Fd���x��� ��$p ȁ3g����r�-�=l7[���ۏ���     �~�����q�n�nnn.  �Ow ��������:Ȗ�Xn٨T�     ������]��nbb"  �Ow �XXX��$ۛ彈ٳ     �l��Yc���  �K� �ɂEK��� ;N$p��b     �fe/�Ƃ��  ���  '���c?{�%yv�-����    �(�V��D�XpwSSS @�� �D��.pϖ�8l���;��ؐ�:    �O�k�Y|�V��� ��%p ȉd�buu5Ȏ�:lo��b���     �~��W�,������  �	� rbff&��� ;
��:�j,�    �S�l�R)8����s��  �K� �.\����+{     �j��Yd���  �M� ���Ӈ��V�dC�@�����c�:ɂ;     ��䆾���;���݌��  �M� �#CCC������J���f�X���~-�V��    �/���7�,������  ��	� rdllL��1'�'�5��j�L�     ����^d���ݜ;w.  �ow �9s�Llll�qR����/p    ��l�ewاT*G777  �7�; @��?>�߿d�I�ɂ;     ���޿���Gg� ��	� r�ҥK����qR��z�     �o�L����y3<<� @� rdbb���f�d�I.�7[�(9�    �'���_oD���ͩS� ��'p ș���(��A6�ԁ��j�F�3��     �`m7���&�D�ٳg ��'p ș��)�{�����nY�    @�X/�EVYp7��� @�� ����L<~�8ȆB�pb���nv�     ���|��]�Ʌ ��'p ș������d�I��v��T+     ��V���jd����J�R  �O� �3�����v;H��<p��עVo��?     �m[��h�Z�U��  �A� �3��tdd$��쮚��I��v+�p�t     @����E�%k����T  �w �����g��     ^�^�D�Yp?����  � p ȡ���XYY	��\�2�h     �5��  ��  �����޽{A�ub�     ���l�N�Y&p?�B��N�
  �A� �CKKKAv$G�f�y"�V�ވ��ZL�     d�zy/��vd���hFFF ��� ������O�^��$���NE�    @f���E�	܏���� @~� rj||<�����+�'��m����ٳ     Y�.pϝ���   ?�  9u��Y�{F���{u�     �U�l����[XX  �C� �S.\��w҇����l��t���     �i{�ß,���w �|�  �.]���y�~�ћ�vlU����X     @���f{�=a��h���N��  �M� �S���V��['����    ��Y/��&�N �|� ����X��� �:q�^�.�{s3     Y�����5�Gs���   _�  9v���{t��͕m��    ȖV��sgnn.  ��; @�%�G��։Cw�v���852     �k�{�l�#��o�P(���R  �/w ��v�Z��w�ҭS����S#��     ��uR�����K�  ���  �&&&���f3H�d�$�i�Ov�fe{7��
�    Ȇd�������d  �?w ������ ݒcw��8�_s�O�n     ���zy/��������  �#p ȹ���{t"p��ۏZ���     ����~4��EZ��ۻx�b  �?w ��[\\�����֩c���n,��
     H�~y��X,���
���P  �#p ȹ+W�į�� �:u�N��    �v�;��������h  �Ow ��:�988ҫs���x    @[�����ӧ �|� �������W���h4[1P�*     �S�E���``@����� �|� ������\�ޭv;Vw�175     �F�;������]�t)  �'�� ��/ƽ{����䓥+�w     �ke��B��v��EN�:  �O�  ���b
�h��A:u�ོ�?�7     ��U�{�  ��S3  Q,ctt4����tJ�u�?BX۩D�Պ�_~     H��A=v�k�/�o��ٳ @~�� ����)�{�%�q6��u�VlV�1=a    �tY��WH�ogaa!  �/�� 8t�x��i�^�ѻ�{be�,p     uVv*�O�1~���b  �_w  ]�z5���?��ɣ��v9n/�     H��>
ܓ!�B�������  �%p ��ٳg�X,F��
ҩ�ϖ&�{��vX     5j�fl��G��䝿�LLL  ��3  s�ԩ���	ҩ���F������x     @<��9g���3==  �O�  �M��.pO�N��m�
�    H��[��'��s�ҥ   �|r �o�~ҩ���[����     i�|[��7�B!fff �|�� ���r�J����{�N�>|/o�F�ՊR�     �K��A��k�O�lxx8���  �=�� �������a��_�~�t��v�ݑ_���_we�sS     ��lk7������;w.  �'g  ~fjj*����t*�J�h4:��?���    �sϷ��o�lii)  �'g  ~faaA��b�񻣁���_��B     @/=߶��GW�\	  �� ��y����C�N�>~o��Q�7bx�     ��ʋ[u?�����!��  8�S!  ?399��p�]�T���n�Wq.M�	     ��[������M  ��O�  ����ӱ���O7��6w�     ��3�{.���  $|z �%sss���J�އ_     ��v;Vw+�o�7�z�j  @B� �K�]�_|�E�>��w����b|x(     ��Vw*�h�����,��cll,   !p �%�ϟ�b��V����[O�>�܉�     ��y��2*p�ӧO  ��� �W������� }�Ƚ�ht��H�@�    �m�;��G�7�p�B  �_	� x�d�]��N�ܟm�     tS�ٌ��^��B�еZ���ի  ��3  ������ }����������FlV�qf|4     ��o���jG���Y�T����  ���	 �WZ\\<\i��u�:�'+�w     �ey��(������  ��� �W*���r�?��Y֭����v�^<     �O�v�	���  O� �k����S�[���N%��f�J     ��S���_~����ͮ\�  ���  �֥K����ҥ[��f�϶v�⹩     �Nz�ٟ��	���%/
���  �=�;  �u�������v;H�B��R)��f��'�w     :N��O���  �H� �k���HT�� ]�7���oG�     �F�����W�כ��	  �Gw  �hzz:=z�K��j���>Ճzl���쩱     �Nx���>}M6��'/��j�/_  �Gw  �hiiI��B�\{y��#p    �c�;t����zI����  ���  �����㷿�m��t9%��ŗny��\�     �	϶�y422�b1  �	� x��8<<���Azt3p_ݭD�ь�R     �IڬT�R�G�������  ^E� �/J�>ң��{�ޟ��_�=     p��l��z{B��zW�^  x�;  �������)�JQ(��nx��#p    ��=������5Y�|Ǳ��  �*>E ��nܸ���o�S�v�՗�����^ɂ{��?98    �I8h4c}w/���W;u�T  ��� �E�b1��ǣ\.�����Vo���^�L�     ��d�����:�k��/���  x�;  o%94~��wAzt{�%Yq�    pR����Yo��ׯ  ��� ��r��5�{�t�0�xc;>�<     p\�v;�m�F?
^��ڟ;w.  �u�  ���/F�X�V��C����^��bl�A    ��Y/��~��L��j���  o"p �%ǭ�� �P(��t˓͝�qa:     �8�n��z{B��jKKK  o"p �-,,�S$�ۓȽ^�w��|��%p    �؞llG���K�Yq���  �7� ��n޼_~�e��q�����͝�7�1X*     ��J� 6*��g����5���  ��'i  ������1��h�����f��6w���T     ��x�����CCC��Ξ=  �K�  ə3gbuu5H�^<o�����    �w�h}+�����.^�  �K�  Irx��G/���[�l��T,     �~���{���/+
q���  �_"p �Hnݺ����t�E�~�h��v9��L     ���h�����/���  �̧F  �d||�� Y�Ղ�K�N�cp����������    �#{��yЋ������	  xw  �lzz:�<y�Cr$�zྺ����a`     o��L^ݍ~����/�r�J  ��� pd�/_��Hr$�V�]�=��X�݋���     ���dc'��v��������ii)  �m� 8�7n���v����W+0�6�     ��Gۑ��_6>>�b1  �m� 8�dydtt4������ա�ǵ��立     ���nǳ����/���  x[w  ����\ܿ?�^����جT���h     ��<�܉z�y p�{�  ��  ��[�n	�S"yҳT*E�_$+�w     ~���ȋ^ӤU����L  ��� �Nb`` �F�{�L�Z������Vܽ4     �:�v;o�D
����ٳ  G!p ��%ɕ�����5�^j��kqjd8     �UVv*Q��c0G���+W�  �� �w�$���˃y��~{�|     ��<Zߎ����ڵk  G!p ��ݾ};~���>-Jo�4p_�    �z�7�"/���x��N�:�$  ��'H  ����`���G�\z+�wQ(z���T�zP�ѡ�     ���QދJ�y!p�����  ��� p,��7������j����IT�pm3n��     ��V7#Oz��j�$�<�n�
  8*�;  �r���{J$+��?��    xُ�ۑɝ�X,/�J����
  8*�;  �2==}x�����hZ�rfe���A�[�    �������8/���\�  ��;  ǖ(�={�V���3�w�     $�mF�?�z�j  ��� pl׮]��@����;     ���v���y2d��o
�B\�r%  �]� 8�[�n������X<00�F�'��zy/v��19:     ����r��{s���?����b�  �.�  [r���������u�^��W6���      ��l�=��$�ᅅ��  �w�5  'biiI��Iྷ�׳����M�;    @ε��x�����z��ݼy3  �]	� 8�oߎ/��2��v�;I��K�{��Y�ƙ��      ��n��A�y"p�I�]���D  ��� p"���bpp0���u���ae#�\��(    @^=\��z{"������	  8�;  'fvv6?~�N�T:�i6{�����F|$p    ȥF��7�#o,���ƍ  �!p �ļ��{�HVb��j�~���A��Vbzb<     ȗ'��h�"O
���+���g��` ��� pb�^���o��V��i��{�'~X��    ���խțdx&	��8}�t��  ��� pb�����Tlll���{������ʂ�>    @���x��y���|Z\�x1  ��  ��d�]��[��ý�K��A=V��q~j"     ȇG����+�###���~  �q	� 8Q|�A�����v�������~��_"|��!p    ȑV7#��0<��N��f ��� p�crr2�����I���j��׶�]��B!     �o�z#�wʑ7�BA���[\\  8	w  N��˗�����I��ܓ/3�n�����    @KFOZ�������s�N  �I� p�>���{���9����w    �x��y��{|�������X  �I� p����xT*��7�rP���F3�J    @��ۏ��^�Qv���  pR�  t�ŋ㫯�
z�X,���@4���u4[�x�����     �)���a��ܹ  pR�  t�ݻw�=��{�'��|]�    Ч��v���yT*�bpp0�nhh(N�>  pR�  t����᳜���Ao$�J��뿌Xۭ��^5N��     ���v9��G��_�p�B  �I� �1q����7�tX���_Y     �˃��ȫa�����?  �$	� �>�@��Cɂ{Z$_p|ty>
�B     ��f<^ߎ�J^�ͻ������  8Iw  :&9h&��z=�O��Z�'����A��Rb�vp�L���D     ��oE�Պ���133  p��  t���\���Ao�%pO�_^�    ����W��O�T���u�V  �I� �Q�o���P�S.�#�n����C�    �u��Z��V"���G��XXX  8i�  :��ŋ100�F#�4؛�V<\ۊ�    �l{��������H����{?  �!p ��fff�ٳgA�%O�
�h�ۑ���     }����ȳa�q���  �N� �q7o���Prd��ߏ4X�.��~-&F�    �*����"��a����b1�\�  �	w  :.Y���o~�V+辡�����q��\     �MV6"ϒ�{����ӧ#w  ��;  �8ϝ;���A��mE�����.^���     ��V<Zߎ<���v�Z  @�� �7n�{$m��J� V��q~j"     Ȗ׷��lF�����͛  �"p �+n߾���o��nݕ,�F�^�������     ��lDލ��F�MMM~�   �"p �+�C�����NU��pm+>�7bx�I     �b�Z;|�3ϒA�R�y���  ��& �knݺ%p���r9=_:4[�x���/�     ِ�Ιwɽ=�
�B���{  �$p �kn޼��y4�͠��xp��ٚ�     #Z�v|��y7::yv����W{ ���  tMr𜙙��ϟݕ<�:00�F#�b{�+;嘝<     �ۏk[Q�����+#9_pOƌ  ���  t��۷�=2<<���=����    ����ȻdLfpp0�*2�r�J  @�	� ��ׯ�o~�ԅ�y���T*�H���������G    ��ک�be�y7::y6==}� @��H  ����Ǔ'O��J�Ӧ�jŃ��xa6     H�/�d�����  ��;  ]�O��O�H�MM�UZ�V�ɷ���     )�j����� ��R).^�  �w  �nii�0����Aw%�2{{{�&�{�çmgO�
     ����V��Ȼd@fhh(�jff&  �[�  ����\���Aw�.pO|�lU�    �B^^^����۷  �E� @O|���H�4z���֗bx�Q     �b�Z;|��|�R)  �E= @O\�p��)σ���{���P(D�ݎ4i���`e#�_�     ���k�����Wɫ�  �Mw  zfqq1<xtW����G�|�lU�    ��v;�_��p8&�/�vï~��  �n� �3~�a|����[�w�3�iܷ�����=}*     譇k[Q�7��^Gͣ������	  �&�;  =3==}[W�ՠ{Ҽ2����    z���������W���  �&p ������K3i\����֗bx�U     ze�Z;|q����<J�K�s�N  @��F  詏>�H��e�A:�����#m��v�_^�ۋ�    �����Z�BrS�k�>44�Ν  �6�;  =555ccc���tOr�Oc�����J��0{��     �Uo6���F�BrO/��G�+�  �w  z����q�޽�{Ҽ6S��㍝X:w:     �+q�h/���F^}��  � p ��>����ꫯ��n�1<<|�8�j�"��z�,p    �o��?�k���}OLL  �� ���ӧO���V�=I�^�V#��o��V�S����     ��m��N���Ť�E�N�v�Z  @�� H���?~���ݓ���5pO|�t%�ύK    @w|�t5�I^���B|��  �"p  �ܹ�����V+莴��<Xވ�./��?�     t�n�v���O��OMM����<  ���(  ��<�y���x��Y����Q*���lF5Z����z�Y<     tַ�ע�n?�k��� @/	� H��?�8��_�%�dŽR�DZ}�d%n/�>�
    @gԛ�x���$���I���\�  �Kw  Rcaa!����V�ݑ���R;��;�t�t     �I�~�H�k��266y4??  �kw  R�ҥK���ݑ��U�z�,p    �o��?���y'ܽ{7  ���  ��'�|�}�]����F�^�GZ=�ڍ�J5����e    @'=�܉���U�Q����3g�  ��� �T����S�N���n���:́{��+�n\
     N�7��_���/��|�r  @���8  �w���������;��=��A������B�#    �II�۟m��>�ccc�Gw��  Hu  �������h�ZA�%�{�5���^^�;��    ����h���ύ��F�LMM���P  @� H�b�333���t^��;9ZD�}�d%n/�F�P     ���lƃՍ�ey�oݺ  �w  R飏>����#9֧=p�����v,��
     ����F���熇��a�$���v�Z  @Z� H��/���`�����FFFb{{;��ޓ�;    �1������Z𲱱�ț����.�  ��  �V�߿?輿.ҴZ�H���Xۭ���x     �n~\ߎ�j-xY��B�w��  H�;  ���'�ܻ$9`'+�{{{�v_>Z�����     ��|�t5xY2����dhh(fff  �D� @jMMMũS��\.�7::��������e����     �h��ˇ/e򲼭�'.]�  �6w  R�ƍ��?�1�$pςv��/���q1     8�{OV�W�c�~���  ��� �j�a������f:�T*>Ezppi��嵸{y>F��    �m�Tk�lk7x���122  �6j  R-	�gggcyy9�d�=�{�Վo����Ks    �����A��HB�d&On߾  �Fw  R��O?��>�,�$p��ގ,���J�Y<�b     �fՃz����Z��ۓ��ƍ  i$p  ������j�t���p��h�Z�v�z#�/�����     �;~�-����}qq1   ��  dµk��/�:/��	*�Jd����Ǎ��(
    ��՛����z�jɚy2 �'}�Q  @Z	� ȄO?�4�ݻ��e��R�^�?�Gk[qi�L     �j~�~��jy[o�������  ��� �	���133���Ag%�{�|�xY�    ��V;�y�����x���۷  �L� @f$+�}�Y�Y�b��)�Z�Y��[��[�qa��    �?�am3*�z�zY~9�R�׮]  H3�;  �1??###���tVr��J������    ��~j��M�{x2��������  ��  d�����/�:+9�ommEV<�؎����	     ^x����j�zccc�'}�Q  @�	� ȔO?�4�ݻ�V+蜡���gJ��fdŗ����s�r     �½'+���)p���8� ��� �)���133���Ag%+��r9�������|�    @�m��by;;7�^8|ɋ;w�  d�� ��IV�?�쳠���7[���x9>��     y��cC1�d||<�"y��ڵk  Y p  s���cdd$�����I�
�h�ۑ�>[�;Kblh0     �j{o?o�o666y����b1   �  dҍ7�O�S�9ɡ;�ܫ�jdE�Վ�/�'W     ���G�35^���K�i^|���  Y!p  �>�����/��j����d)pO|�l5~�t!��q    ȟ��~<Z��l||�0rσ����  �
�  �444333���tN�k�V�{�]�    ���ӣe��o!	������  Y"p  �>�����ς�)�J1<<�Z-���+q{a֊;    �+����qm+x�d�=y�4�;����  �D� @f������H��������������%+�    @~|�x%Z��Q�zi�X�<XXX���+  �C� @�ݸq#���?����5_?]�ۋ�c�T
    �~W�����������G^|���  Y#p  �����9���h[�阁������ȒZ��<]�_-]    �~�������R^�����  ��;  �688�����ɓ�s����//ǭ��(y~   ���ޝ>�Yh�>��-�؀1�;lll�l�Kg��d:==�n*5U���n:@��8x��]�*˖dk�۷�3�tX$Y����qT��*��`]��9/(�����>/��ͩ���?�y�  @%� P�������]X>E�>44�JS�����'}(     eu���L�Xo�����T��e�'�x"  P��  T����tvv����ayK�������J�)Vܷ?�&u�V�   ����ʩ�7���.�@� @%� P
�v��|�Oq�_�"(��-.w��    �l������������]ʮ��f��  *�� �Rعsg>���LLL��Q��{����e]�w    �TƧ���/@[[[���u����  �Tw  Jc˖-9r�HXŲM]]]���SiF�'r�ʍl[o�    (����f��l�j܋���{.  P��  ����?�cǎe�S�˦XqN%��lYכښ�     T�"l?y�z������X5oooOwww  ��	� (��p�xv���?,�J�G���Vܷ��    @�;r�j&����W5���~��  @�� P*�/~�<���R[[[�+�8?���Xq    *���T�Xo_�bټ슅�͛7  *�� �R���Igggn߾�^MMMZZZ2::�J426�׳��5    �T�/]ͤ��y����p)�'�x"  Pw  Jg׮]�����hmm����P��oYד���     T���9i�}A�a���)�G  ��  ��Ν;���gbb",�b����6333�D�����ky�ч    Pi��x%Sz>��TC�nݺ466  �@� @)mٲ%G�	K�X�)"�J^q���@���MC}]     *���DN]�毾�>���)��{.  Pw  J���ϱc�*ve|�kkk���}|j:G.]ɮ�    �R������Ά��������tww  �B� @)544�=�����^��^[[[� 8z�jv<�P���    ����z3,L5�O?�t  �L�  �ց�_�",���֌���RMLM����ٳ�     �t�����>MMM)�b�g��� �2� PZ===s�r�����Vс{�X���|dmZ    �R�˹�Caa�;��۲eK  �l�  �ڮ]�������ܜ���LOO�RMM�����o�     �T��d�z�������jjj�{��  @�� (�'�|2�|�I&&&��kmm����������1     +����\�q+,Lcc��W��_�>���  �ǿr (��y�#G������V����L�p�r�o},     +͗���}���w��  @	� (�����رc���	K���infjj*���������t�6    `��6<����yP��www�} @	� (�"�޸qcΜ9�^��~�Ve?�;;;�C�rpǦ     �_�W��444��jjj�o߾  @Y	� �
/��bΞ=;2��Z[[+>p/��v3?ذ.��Z    ���Wn���+�z{KKK֭[  (+�;  U���z�\�|9,���ƹ%����T���_���kOm    ������8eܟy�  @�	� �Ŋ�����Yq_mmmJ��pchn顮r_~     +[�����ݰp��ͩ�/oS��lݺ5  Pf��=  �'===����͛7��*K�^����yg��     <3�����H����;v8� ���  T��>��կ��*�p�՘���T��Gs���l\�*     �۱�k�S�����.O?�t  ���  T��{,����s�NXZŊ{�B�⾡�;�55    �_&��s�╰8����զM�R[[  (;�;  U��g��o~󛰴����7o�F�&r��Zv>�6     ��.\���Y�2�����d�޽ �j p ��<��S���2>�ץT__���挍����kW����M    ��+�7N\�S��K�e������1  P�  T��۷�СCai�e	��'��޳�     ,�/�dfv6,N��^[[��z���  �B� @U���Çgz�S�K��3[�K����d��k��d    X>7������a�:::RV===�^� ��L� @U*V\�x≜<y2,��	���֌����gf��������     ,�b��ū��OKKK�j߾} �j"p �j8p �N�*���JQ<[���p��`v>�6=�    Xjn���[�a�ʼ�^���Y�&  PM�  T����<��ùt�RX:��X˙��J�����y�m    XJ���W筷߫2�{��	  T�;  U�^�����3,����ܺu+eqyh8�7o��U�    X*���֝��x��JCCCʨ��6n�  �6w  �ڪU���ӓ7n��S<�Z����Y����=;SSS    �{55=�?\��M��۟z�  @5� P�^|����K���>MMMOY����+�ٲ�'     ���+�;1�$)Wʨ8g߱cG  �	� �z�֭�[xK��T(S�^���<�fU��j    �Xw&&s��Z�7mmm��-�y��͛K�� ��� ��ڿ���1,����fvv6eQ\:�x%�l\    ��:t�r��g½)�kʨ۟{�  @�� ��ڴi������hX�|���w����y]Oښ    �P��w�wu0ܛ����3�2�� @�� �������{/,�2~h`zf&�����;6    `�~�w�T/_>(e^o߳gO  ��	� ��mݺ5}�Q�޽�FKK�܊���t�����l[ߛ���y�    ,���n���r��<(e�7nܘ�F/� P��  �<��s�����)V�o߾�������ճ;RSS    ��353�/���{���T��8o޿  ��	� �?عsg>��3+�K��������ȝ��|=�֯	    ��9|�JF�'ý+�z{}��  ��  ��ݻw�w��]XsK:)�/����5����    �#c�9�5ܻb�V)���z���  � �/<�������3>>�Fq�088����ʡs����G    �m>?۟��p����RWW��y�G��b   �;  |�]�v�O>	K��o޼����]�뿚-�{���    �����p.ܸ�FgggʦXo?p�@  �#p �o�{��|��WVܗHq8_�ꌌ��lffg�ɩ�y�m    �����ߟ�K���>---)���ק�و
  ���  �œO>�/��",����R�[`ʆ��     �щ����FWWW�h���  �D�  �b�޽���399�]cc�����D���������    `bj:__��F�Rh1�R6�֭�{  ��;  |���ڹ����*,���������s���`ú     |q�?�S�aix]]]ʤ��8  ��	� �;�۷/����T�wE�~�����Φ�������!    @��9z7���s��A���L٬Y�f��  �sw  �Ŋ�����"w�]�FS�쌌�����g���Kyi��    ��gg.�v��A���OKKK�f���  ���  �G�<���ǭ�/�����+7�m]o�vY�   �jt���\�U�3����+e���[ʟ  ���  �G��e˖;v,ܻ��ƹ�����է}����s��    @���W���*�S��?�a  �o&p �yx�r���LOO�{W\Fܸq#eucx4'�g��k    T�C�rgb2,������եLV�Z����   �L�  �P__�'�xb.r��������MY}~�R6�v���!    @�����������J�8p   ��� �<�������jjj�"��������t~�w1wl
    P~�������z<��LKKK��z;  |?�;  �Sccc�mۖ�G��{���Q���p��`�X�:��.��    �'���ȵۣai�q���^  ���  � Ŋ�ɓ'355�M��kbb"eV�6�������    (���|yn ,�b(�L֬Y�իW  �nw  X�����ر#_�u�w��č7Rf�w��������p    ����̥�OEYjmmm���K�8p   ��� ��߿?'N�(����P\Pfvv6e��������jm    P�n����`Xz]]])�u�֕�g ��"p �*Vܟz�|��������E�###)����|r�|�|f[    �r(��>��^CCCZZZR&/��B  ��� �"�ݻ7����d�7�����C�9{mpn�    �|G/]��ѻa���e��#�̍�   �#p �E(Vܟ}��|��'��K<���K�}z�b^ՙ�z�   @%������W��Y����y�� �¨*  `�v�ڕC�UE���:::���xwb2_�Ⱦ�    T���.fjz&,�"n/Ff����y  �O�  �`߾}���½immM}}}���Rv���eӚ����-    T�����XeZo/B����  X�;  ܃;v����}�ܹ�M��~��͔���l>>}!���>�4-    P9�ff�Yߥ�<�1���ƔŦM�J��  ��"p �{T����?�s�7���������hN\����    �89��aytuu�,�������  X8�;  ܣ͛7�O>���HX��ֶ����=~q�?��v���!    ��74z7�������0��^[�lI}�,  ÿ� `	����?���T���r��쬚�}bj*����W�|"    ��V��~�w133΀�K������  `q�  �{�ttt����a񊅞��挍����~3��-�    +ױ��v{4,�����3��عs�ܫ�  ��� `����������{S\bTK�^����<�՞��   �J4:>�C���)^�,K^__�ݻw  X<  ,����g�������:w055�jpwb2�?s1/l{<    �������	˧���駟��v  �7w  XB�/����Ά�+V�o޼�jq��<�fu^U�K    (�SWnd`h8,�b����1eP�E�  ��;  ,��kצ��7׮]���ޞ��������N��}��4��    x����8��WWWW�b���  ��  �ث�������W��/^�|k[[[FFFR-F�'�����ۼ!    ����鋙��˧��an��ZZZ�cǎ   �N�  K���;6l������uvvVU�^8�-{WemW{    ������0x+,�2���߿?  ��� �2x���������LX�b����9ccc�����N��O�<��ښ     ����t>��WMMM:::RE�_�   KC�  ˠ��1۶m˱c������n�ˡ�y��    ���]���TX^�+����)�_|1  ��� �2)�O�>���ɰ8���sK���;<|�r��NO{k    �����휽v3,�b��z����  X:w  X&����ݻ�駟��+V|nܸ�j23;��?��zv��T    `�MM��Ӿ�a����ύ�T����<x0  ��� �2*����:w�����֖���LOO�����#����    X~_�����DX~eYoߴi��K�  ��� �2+�[���1���a������Ƚ�|y�?z����    `�\�=��W��%����%��ͩtuuuٿ  ��'p �e�q��tvv�֭[aq�����Uۇf�����sy{����    Xz�9�G�.�H����ݝ2xꩧR_/� ���_�  p����������8���ioo���p�M�u|�Zv<�6    �����@n�˯��1����t�ϱ{��   �C�NU�  ��IDAT�  �Aooo֭[�˗/��)V�1p/|�w)�;��Z���   �JRL����ٳ'  ��� �}��k��o��o<s�H�S�mmmM����ɇ����۵#��5    ����L>:uޙ�}RWW7�Rg�+~�m۶  X>w  �O�C�M�6���/,N��^��{����x%O?�.    �����K�}w<��z{MMex���  ,/�;  �G̹s�2==���1���K5��|^Ց���     �704�SWn���Ë�J�z��_�>  ��� �}T�O=�T:�����}ff6�9q.�����V��    <(�������p�tuu���6���_  ���  p��۷/Ǐ����o���e��FC�w�չ����H    ������ܙ��O�W�G}4  ���  �b����?��ð8Ŋ����S�_��GVw�.�)    �o�쵛��)������S�s�^x!  ��Q�A  @�ڹsg��⋌����kmmM]]]���S�fgg����_�>�����    �����puww��mݺ5���  ��;  < ̯~���p555s+�7oV�����x~�w1�o},    ����ԅ�OU�hƃR��466����ū�  ��#p �dÆY�vm�^����=�n����L���ky��+���
    ��N]��K7o�����{��Im��4 �~� ���o��?�yUGڋU\(�����})����_�>���   �7���g�����Ԕ���T�����ر#  ����  ��x�u�֭9~�xX����gvv6����d>9}!wl
    �犳�ߝ<����p�Z�*����&/��R  ��O�  Xq@~�̙LLL������[q/"�jv��`����5�}a    K����\�5���ƴ�����[�.k֬	  p�	� �����������������HU��>:u>k�����     �}w,_��_�����  �`� `ؾ}{����ܾ};,L��^,�{5���G'�絧6    ����l~s�\�gf�����0��f%{ꩧ���  ��� �
��(��n�/�/F��>::Z���7�r��Z�?��\    �ۗ�28z7����^���>�l  �G�  +Dooo}��\�p!,L}}���Y߅��jϪ��    @5α�k��+�j;::R����  ��� �
����g?�Y�����+��dzf6���O��L]mm    ���ON�w'��K�F����^�:�=�X  �K�  +Hccc�y�|��aa���>::�jw��X>뻘緸�   ��|t�B�NL������kjj��+�  x��  ��<��s9~�x�ܹ�Xq��������l��
    T�c��rq�Vx0����"�J���Wt�  e"p ���_ί~���0imm����g�=;���    (��U�/�����.����T����/  X�  �mذ!����~�zX�b�]��o�'����y����    �ezf6�9q�_�;�J_o߻wojkk  �w  X��x�����?2;;毱�1---�{�nH����+���u   �2�����u������H�jkkˎ;  �w  X�:::�e˖�<y2,L�$p��/��g]wGz;�    erq�VN]��J_o?x�`  ��E�  +��/���g�frr2̟�?73;����O��LC}]    ��NL棓�ÃS[[����T����g�ڵ  V�;  �`����������)�������x>>}!/m<    P�fgg���3>5�b��8ǮD��]��   +��  V�;v��/����p�����477gll,���+7�pwG�x�'    PɎ\��˷��>HE ^�T��۷ϝ#  +��  *�o��w�}wn���+.W��S���ٞ�7    T�#wr����`篕����ؘ�{�  X��  Pz{{����̙3a��w+�njz&;��wmOmmM    ���[�=q.33�@�"l���N%����K/�T�q>  T�;  T��_=?��O399毸d�|ٚ�t}x4_��ϳ�	    T��O_�����*�]+5_�vm}��   +��  *DqY��/�׿�ufg��WSSSZZZr����'�p9������    �'/_��k7ÃU�UwuU�b���k  V6�;  T��[��СC�W�		���oO��O��L[Sc    `%�9z7�?��U�VU�z�3�<��F�  ��	� �¼��[�ۿ����̄�).,Z[[s�Ν�'�S��Ѿ���m���)    �orz:�;�ig�\]]]Ů������  ��'p �
��ё;v�ȑ#a��w��_�~{4_���s�    �D�;y>#c���[�zujjjR�^}��   �A�  ���������X��������ett4��#��dmW{��    �$G���[������`�D7n��� �� p �
T[[;�6�_�*��W�gggß����j��_�   �����h�<�V�J]o������  T�;  T�6d����S,+�###��MNO���}y�����    <HS�������X�2+q�����΍�   �C�  �7��_��_gzz:�O��>::j�����O�.f���    Jqv����+C��^����[�  �,w  �`���ٻwo>��0?�s�����D����h��    �×�f`���J���8w�Zi����^{-  @�� @�۵kW�9����0?�jO������>:u>��[���    ����ɡ���Q���۶m��0  � @)���y��w��T[[����ܺu+������h_�yvG��    ����T~{�s����)mmm�4���o߾   �I�  %��ۛ�7��ٳa~��}xx8333�/ݺ3��N����    ˭�ڋ����dX9zzzRijjj��/��   �I�  %��(?��O39�h>���>44�ٙ��y��=�֯	    ,�C.g`h8����iiiI�Y�vm}��   �K�  %Q�����|��o߾m��;|z�Bz:����    X�7o��ūaeY�zu*MqN�ꫯ  �lw  (�;v����߯x����+7o��lzf6�r�t~�gg��		   ����oO����lX9Z[[+r��駟NSSS  �ʦN  ��y뭷���V�穣�#��Ù��
߬�d|�h_�xz�܇    `)L�����g2>�ln����I�iooϮ]�  T>�;  �Ll��?ȡC���+�����\�~=|����|q�?{6=    X
�;y!��w����ٙ���T�����_  Pw  (��>}}}	߯��mn�}||<|��/\����<�fu    �^�t5��+K��^]y�۶m�2  �A�  %���8���������ˏ+W���������Ҝ���    �b\�W���S����ե�477ύ�   �!p ��*Vv�՚cǎ��W\������]O"�陙�����ɞ�ij�'%    3:>�O����lXY���W�_{�   �F  �{��s���ܹs'|�U�V	�硸�|�h_�xz�ܓ�    0�x����d|r*�<�hJmmm*ɦM��f͚   �"p �+.#�|����̬E����А��������604�/��gϦG    ��ѩ10�g�����$���s#/  @�� ��֮];�b����_�������.gu{K_�:    �]�^����n�����'�楗^���y  `~�  P^{�\�t)������ե��+CCC����Ĺt�����%    �M.��saejnnN[[[*ɣ�>:�  ���  �@�b��������+�����t�nS�3���O�'{v�����    ����|x�\f���b����������_  P^�  �Ś͆r���jjj��ݝ7n��W\R��/o<�u�w    ��ټ�L�'�����ޞ���T�^xa.r  �˿� �����[��O�����݊��۷o�]��@�����<��    @��28r7�L�X��իSI֭[��<  @�	� ������W^�����7|�U�V��իa~�p�rV����5�   @u;r�j�������+�uuuy��W  ���  �̦M���C�ʕ+ỵ�����9ccca~~{�l�Z����%    T�?����U��tww�Rk����Kccc  ��� @z����,����+�a~��g��_��_�ٙ�r   T��w����3������Y��s�b�R��m�  T�  T�b��������w+~Wmmm�3:>���T~�k[�kk   @u���ο9=�_V����tuu�Rk��z  ��!p �*�s��=z47n�߭X�s�Nfgg����o���+;�    �733�����[pge��驨u�ݻw���5  @�� @{�����<333��O��FCCCa��]��C�yf��    Pn����˷�����Ғ���T������?  P]�  PŊ՛�{���O?߭�H���T��/�����)�֮    �t��՜�V����T�be�G?�Q  ��#p �*W<���ח7n�oW\��Z�*׮]����"�ގ�    P.�7o狳�a�+F<S)v�ڕ���   �G�  �w����s��ߣX�onn���X��陙�w�t�yvGښ*�   ��v��X><~6���ae�����Օ��bwww�y�   �I�  �E�/��B����݊K��~�Tuwbr.r{�����   ��6>9����ebj:�|Źf]]]*A���  ���  ��}���8q"�/_߮��a�Y����0�#w��3y��'RSS    *���l��h_F����W�ivuu�����{M  �^w  ��y���������d�v�󸣣����	s��P�8۟=�	    ��S�s��h�������Z��   �M�  �?Œ�+��������l�f��E�>88�����ܘm��   ��r��@�\u.V)���*f���.?�я   p  �̦M��裏���uttddd$a�>9}!�-�Y��    *���C9t�r�555���I�8p�@   p  ��[o�����g�nժU�r�JX�����������t�4   ��mp�n~{�\��+�ū����G�O<  ���  ����y��������577�=�{�Ν�p�S�y��鼽k[��y
   �Rݙ��{�Ogjf&T�����������W^	  �)  �o�裏f���9}�t�v�W��ݻw3;;nh�n�;җ7�ޚښ�    ��L#�O���d����sC&���_���  ��_  ��z��W���?p�͊%����ܺu+,Ε��|x�l�x<5"w   �cfv6�;����+I��d{{{*�ƍ��V   �#�;  𭊅���~;��������Օ���LMM��9{m0mM����,   ��⣓�304*K��^	�����  ���  �w*.Cv�ؑ�G��oV��www����a�_��֦��|dm    x�>?s)}WCe)^�ljj�JW�����ks#+   ���  �^/��R.^���akMߦ��-###��Y�Ŵ55���    �`���#����R��W�N%غuk֬Y  �o"p  �����/~���̄oV\dvv6,N���ؙ���֬�l    �ץ�����b�<===����J��ښ���  ��� �y�����ݻ��矇o���0��[���M��佯O���;���    ��w���3*PSS���d%x�7  �]�  ���ݻ7}}}
߬��+������
�7>5���d�yvg���
   �܆���ޑә���c%Z�fM*�~���1  ��   �w������df�E�7�����իs���poF�&�"�?�=�u�   `y�ON�ç36i���x���� {��	  ���  ��֖W^y%��^�f---imm͝;w½)����Ѿ�������   ��553��������Py���jժ�tuuuy��7  0w  `��lْ�'O��ŋ�+�ccc�����[����غ1    ,��������\����7��+������ύ�   ̇�  X��������ܽ{7��b��xr��͛�ޝ�����<���    �4>�7n��T�ŋ�+݆�y��   ̗�  X�b���λ�;���_������h&&&½��l�\����    po�ȉ��2���̭��t���y�W  �w  `ъ�ݻw�/��l��չ|�rX�;y.-�yxUg    X����9tޙU%[�jU����o�97�  �w  ��<��s9w�\�_jjjJ{{{FFF½���Ϳ>�7�ޚ�]� ��ٻ�/9�3��w眣��X�!
!$�P ���?p�Ú��0��$�s@����\������P���:��>�խ�9����} ��|:4��,_I������ʅ�   ߖ�  �iO?�t���G����%�8�����f��������������Z_    |3�����";7,_�������-���   �.�  �M�����<>��do��c6��_~r&����h��    ����d�{�|d���嬡�!jjj"������ݻ  ��  �b�ڵ�~���p�B�����cbb"�����1�J�[G?���*   ��665�;�L&X��A�d�|��#�De��:  ��  �&�������Bn�Qkkk���Ɯ��f|z6���I�U��   ����T�u�lnX �[�'����ƍ�[n	  ����  �7���{��K/��l6�����hll����`��LN�[��ƞ;7GyYi    �T:~�ə����������b>�����z(   n��  �W---q�������555�&ܧ�&fͧ�c�5ۻ���%%   P�R�Lnr���L�����Dggg�d�ɓO>   �A�  ̻��;.^���%�Q�*����`~����{��ǎ;6��  ����f���chb*X�������2�Ur����?  `>� ��o߾�����F*�
����:���c||<�_WG�w�/�C��   �b���ůN\��1gO����"�53�%����   �/w  `A$/�J�W_}5���/K.����"����\�`T���}�   @�����:<�$/��m��9�]�  `>	� ��bŊؼys�:u*�����hkk����`���:5��mMw    �?��������Ԕ���v�����  `~y�  ,�G}4z{{cl�Ԩ�WSSuuu111̿#��&�o^�    ��K�q��0�B�D㭭��϶l���L   �O�  ,�����?�t:���jjj*��l0�~�J.r_בߗ�    7�T����J_P8:;;s[ �UKKK�w�}  ��  ��K&�?�����o���\�W�%U�_�~=����oO]��X��    ��l�`��ܕ�p444��T�U2]��'�  ��"p  �ڵk��n��'O_VWW����/�_&������wl�   �|�`�^�^P��ʢ��=�ٮ]����2   ��  X4�<�H������p�e������f����"r|��X��    ��������LGGGn�c����;���+   ��  XT���G�J���J&3577���P�0��������m����!    ����G�7�.FV�^P���s��U�o߾=   ��  XT���ݻw�k��f���ihh�����$wF:������]�6EW��   X~z����(���������"v��   �A�  ,�U�V�V�~��������EOO���3I�~.vo�5��w"   ��K���N���$nO�<棒��x�'r�K   ��  X��\�z5��*//����N*��_=���m"w    ���܈�N\�LV�^hjjjr��Q��{ߋ���   X,w  `�8p ~�����l�W���199333�M�s��w�m��   ����s��3�lPX��<��񮮮�6N  ��$p  �LEEE�ݻ7~���Ŝ��_���}}}~.l&��_~r&����h��   �|sml"�9v>�q{!jkk˝�棪��x�'  `�	� �%�����sO��O
����2���bdd$XXI���G��ɻ7GSmM    䋡��x���He2Aᩮ�Ν�d���={���4   ��  Xr۷o�+W�D�W�����T���k:7��l�{s4TW   �R��_=�iq{!J򮮮�W��{o���  �R�  ya�������s�������鉹��`aM����NǓw��Օ   �T�'��-q{A������L6V�^[�l	  �����  �����ݷo_��'?s���+��444,�\���\�^W%r   ���L�}�\̈�Vmmm444D>�����{,   ���  �ɴ�x ���௒ˮ����o|z6���L��֨�   �hlj:���lLͦ�����|TRRO=�T�5  ,%�;  �W�n��.]��W����===��f���\&������E�   �������(++�|t�����dy  ��� ���L	�я~db��H.�ZZZbpp0X3�q��S�����P]    eh|2�:v.fR�p�����Ѻu�b���  ��  @�IV�:t(^x��d2��˯$�������l��t.ro��   �ohb*�:z6f���
Y2����=�Q2���G  �|!p  �Rr��k׮x��7cnn.�\kkk����Q2���OƓw�M��   0_���<z6f�����3�����ػwo   ��;  ��֮][�n��G��K.����ڵk��N�㍏NŞ�6Gs]M    ܬ���x���H��^ccc���F�)))�'�x"��u   ��  �k<�@.����>�\�������D�xr��ǧ�m����.    �����x���Hg�AaK&����E>���r��  ��  �{����^��7�)���ӑɘ�fR�x��ĝ��]�   |=�c�މ�ɊۋA����F�I�g�~��  ���  @�K.�8/������$?���v���l:���L��vkt4��  �o���|d�sA�knn�����7�cǎ   �Ww  `YH.]v��o��f�͹ LTWW�~.7n��l:o~r:ߺ)��   �_�:�yܞu�U***r[�Myyy�ݻ7   ��  X6���[�n��G��kii����H����Jg���ѳ��6�;   ��.]�ߞ�(n/"]]]QRR�$y=O<�Dnp  @>�  ��<�/>��joo����`񥳟G�m�+[   ��]�6$n/"�������7��{otvv  @��  �΁�?��?brr2��eYsss����/���9v.ݲ>ִ5   �.��g.ǜ��h$�ѓ���&َ�e˖   X�  ��SZZ�^x!2�L�����ӹ/_&������wl�   9�{���_���ܲ��+�MCCC�ر#   ��;  �,%�2;w�z�%�ioo�����f���K֌�{�|�ۭ�ĭ��   �c���_.�ť��#���+�H^�޽{  `9ɯwV   �����c�֭q��� ���,����ڵk��H>l�ӗ"�����oZ   ���\�ǯť��1���#����Į]����:   ��;  ��=��100��"���6w�6>>,�?��4�S����U   ���?w%��ť��"�]1�|�{ߋ�.C  ��G�  ,{���G155D������L�R�`�����LܿiMnZ   P��ss����HP\�s����;�Y�fM�y�  �	� �e���4:/��Bd2�(v�eZ21���/79��s��Z�>��|h��~O��   ��L6~u�B��ŧ��-*++#�444�Ν;  `��  !��y�����u&�Tknn����`i]�Mr�qǆ(/-   �p$���9~.��Mŧ��6���"�����޽{  `9�  cÆ144~����3���1==SSS�Һ:4�?:��m��
o�  �Lͦ��c�bx��K1*++�����'�f�={�Duuu   ,gn� ��r�����`\�|9�|Eroood2�`i]�1o|t*��ks�VV   �|�O��[G�ƍ陠8uuu�"�|���F{{{   ,ww  ��<����/榹��-����729�x2vߵ9��   X~F?{��퓳��8577GMMM�-[��ƍ  �� ��t����������t�䲭��!nܸ,�d������w��u�u
   |�������1��-�XUUUEkkk�U�V�}��   �B�  ����x�g�^�LƅcKKK������l���fS��ǧ�񭛢��.   ���7r#�=q>ҙlP�JJJ���+�g������;w  @!�  +�Z�{��x�7bnn.�Yr����===E���3�t����x쎍���1   ��u��p��Rd��U�Yr�VQQ�"�q���(--  �B"p  
ښ5kr�y���?D�+//ϭO�C2���g����Ǻ��    ��ɞk��W(rɤ�d�F�H����z*w�  Ph��  
��wߝ��ϝ;�.��������� ?d���W'���䊸{��    ��Ǘ{?���[2�=�ޞO}��hnn  �B$p  ���?���q���(vmmm1;;�T*�]��t&�ݰ:JJJ   X:���?}).^�[rN��Օ���/����rK   *�;  P48�?�|LMME1K.咉S���Vk�Wbbz6ٲ>����   �I��wO������������|�v��\�  P��  @�(//�C��/��L&�Y�V9��n�}��<8o|t:vm�U޶  �b����w����������룱�1�ESSS�ر#   
��r  ��444ľ}��W^)���uuu1==�㦑��7&���'��5�3!   
���T�}�\LΦ*++���3�E2E~�޽  P�  @���z(~���}��������/�ˍ��x��S���M��P   �����:y!f�Ž��ϕ��DWWW��|PVVO?�t.�  (w  �(mٲ%�������Q̒K�������l6䗩�T���xtˆX��   ��;�?���lqB௒�|�ɓ�;wF}}}   �;  P��)����Ŭ��<����ڵkA�Ig��αsq��5�yeG    ��dϵ���O�����/���X�re   �;  P�����?�|LLLD1����]�ݸq#�?sss����1>3�_�*   ��������O�t���/$S����#_lڴ)��  ��� ��VZZ?����?�q���D1kii���٢�9䳣W�bj6ܺ���ݒ    ��d[گO]��Cc_H�	�����$?�\�����  �b$p  �^uuu<x0^z��d2Q��˻������l6�s��193�ݱ1*��   ��fҙx����6V����G���QQQ����>v��   �J�  ����طo_���Ew�����0��w�F��t�ܺ)j+���   ����t�}�|�O�^Ǘ%g�uuu����r�8���   �J�  �_��;v�w�}7���X���Dccc��Yӝ�oL�/����[7F[C~\�  @�J>,��c6��[IP���� >���(/�r   �ͻ"  ���iӦ�q�F��O�b���333�/���l*^��T<�y]��̏�X   �7g�����l�4�%Sғ�%%%K�Rr�婧�ʛI�   KI�  �w�oߞ�^~���(f����l6�_��\���ܚ��׮   �sɆ�/�ƱO��JWWW^LKO�Gy$���   �;  �WڱcG.r���b��D������܅0��K�165n^e��   �,���oN]��Cc_���5jkk��e���{�7֮]   |N�  �O<�����/���H����hii���� �]���عuSTWx�  @qJ��s�|�NN|�$lOμ���͛c˖-  �_��  �'JKK�СC���8����X544���l�������D�z�D�ܺ1Z�~
   ,��}�{'��t*�U***���+���5k����   �L�  �5*++�?�A.rO�RQ����I�|��&ff���N�#���5m�   �����ݙK���|���������Xj��ͱs��   �	�  ��de�����_�l6�(����쌞����,7�L6�=~>��[��t   ��/�~���u����@��VSS���   ���  �H&��ٳ'�x㍘�+�)`eee�Ƚ���h�M��t��ո1=�o�%JKK   
I��ߞ�WG�NKKK���-�ˈ���8p�@^L�  �Ww  �oh͚5������_��wUUUn}���p�|��c�������Q    �ar6�?C�S_'�И�XjIԾw�ި��   �9��   ��w�7n܈�?�8�Uccc�R�������Ň'�񭛢��%*   ����d�{�|.r���LL���Z�%%%��O�G   ���   �����###q���(V�ī�����Ǎ��x��S�����!   `9�pm8>8s92�l��I���������~<�@�   �	�  ��'�|2^z��b�\�uttDoood]&/+3�t��3�}��ضƥ*   ����\|x�7�}��MtvvFee�R�����cӦM  �7#p  ���y�x�bll,�Qyyy��?w����}�p5�����뢼li��  ��2���oN^�ޑ�DKKK���/��ȅ�w�uW   ��	�  ��d���>���'''�UUU�.������������[7F}uU   @>J>����b|z6��������֥~�f͚x��  �oG�  p���=�\.r����b������1>>,?�S��_N�#����-�   �$�p�g.G:��&***���k�_Ftww�Ν;  �oO�  p�����?�A.rO�RQ����r����L��̤���O�Ķ5�����   �Zvn.>���>���JJJray�yq)%���   |7w  �yPWW���_~92�L��򰣣#z{{���/G�����t<|ۺ�(/   X
��}�b���6�����ť���O?�t   ��	�  �I2�i߾}�ꫯF��f���Gggg������\�<]�_|x2�cc4�V   ,����x�ą����6Z[[sC(�R��1�ۗz�<  �r'p  �G�
�ݻw��Ç�2򮪪�����~�z�|%Sܓ�����ǚ��   ��p��p����H�� nN}}}n��RJ&�'�z�<  @!�  ̳[n�%v����^QF�Ʌb*�����`�J�3�α��mMwl_�2JJJ   Bvn.>���>�������V��TVV����   ��	�  ����333��e�L�J��111,oG���&�?tۺ�,/   �O3�t�������m����6*.���駟�}   `~�  ȶm�r���#G�����"��g��vep$^��d�ܺ)jL"  `~�O�{����l*��J��+V��RZZ�w����   `��  �=�����q���(6�%c����7����LN�+GN���ƺ��   ��q~`(~�Jd�ـ�+*++��5<��c��/   ��  `�=��C111�.]�b�L�J.����"��z�Ke2��o�#�۸:�JK   ��t&���|W������%}?�p�^�:   �w  �E�gϞx�Wr�̋M2I+�t
���k�5�;�l��꥝�  ��165����UCCC455-�󓭅۷o�6   C�  �H���/��rE��������6��Pޘ�W���o_�Z��R  �����P��ܕ�w��������cI_�w�۶m   ��  `����Ƴ�>/��B���E�I&k�R�
�L:o=[Vu�=�W�;^   �2ٹ��ūq��Z�ͨ���+V�&�/�M�6�=��   ,,�;  �"J"������8&''�ش���"�����p��:C�S�Ȗ�Q[Y   ����_���S7#9SK���ϥ�v��x��  ��'p  Xdɴ��{.7�}zz:�I2a���+z{{s�;���F��������ʖ�   ��]��\��t:�fuww��ԖʪU�bǎ  ���  ,����������ܓI[�����=���c&��_~r&�����V.��p   �Fvn.�\�'{�̇������Y��'q��]�  ��#p  X"I���$����(&�ĭ�rr`` ����r�J_ޘ�G����
G   �bb&�>y!�ߘ�����ظt�����cϞ=  ��r�  ��jkk��������Yt�{2y���%������;2�9���;�  �����h��R̦3󡮮.��ږ��ɳ���   ,>�;  �K.�I�/��b�E���L&���Aᙘ�����;o鎻nY%%%  @a����6y}r�ߖ6�MUUUtvv.�󛚚b�޽  ���  ����8t�P���ˑN���$Sܓ�}||<(<I��ѥ���o_5�  @aH>���S�b`�{z�Oyyy�X�"JKK���I�~���%{>   w  ������<�L���?�T*�$Y��D�SSSAa��?���x�u���)   X�._��^��t&`�$Q�ʕ+���lI��l�  ,=�;  @I��<x0~���bQRR������Aa�N�㭣gc˪����UQ�  `�Ie2q�BO��0���dr{E��l���˝ˉ�  ���   ϴ���.�~���U�\vuuEooo���p��:�[_���룱�:   X��'�7�.���L�|K΅���� �۟}�Yq;  @��  ����ؿ���?�l6�"Y?�E�^L�w1�1?���$�d�;   ��dϵ8r�jd���[r�D�K!��:$n  �#w  �<���{���^{��b�du����ǜK�������D��x�ֵQU�   �L�����K�3<�ZZZ���iI�����<�L��;�   �'ޥ  䱕+W�SO=���zQE���b2��ڵkA�|}$������GWS}   ����g.�L:���룵�uI�]UU���+++  ��"p  �s�V��'�|2��D�d-u:�������O���O���]�+���$   X��\����8���,��������D��  �)�;  �2�z��صkW���[E�'�3�L��Y�^���W��o�F<�e}�WW   �ktr:~s�bOL,�$,������{���6  ���   �����2rO�T'��'''��p��D��ȉ��-��si֔  ��C�W"��,����X�bE���.��+**rq{mmm   ���   �H�?���_���"������닙���8�ҙ����?z#�۰&����  �X̤��3��ӡр��D�+W�����O��   ˇ�  `�ټys����.��=YW�������J���q��z���÷����   `~���g.����,��|���;*++���3��   ˇ�  `ڰaC�R0�ܳE�6<����ٙ���d��113o||:���{6����~�  �9��#{�L���Ő�����,�s��   ˏ�  `�Z�~}�ٳ'>\4�{�J:��D���=�W'��&>|��h�w)  �]����N_��3����-�����I���3�Duuu   �|�  ��5k��޽{��^+��;��L"���������x�/'��]�+���4w  �o*����/���177�Z[[���yџ�D�Iܞ�%  ���  ���+W�����W^)�໪�*����ڵk.�P����W��o�F<�y]4՚�  �ޘ�ߞ�cS���x������eџ[SS��  ,Sw  ��L4?p�@.r�d2Qjkk�;r�8]��W����׮�������4w  ���|H��Ձ��rod�>$��ihhȝ�,�$n��g��\  �\yG  P :;;s��_}��H��Q���rS�������ȅ����h<tۺh��
   >7:9���>4>���3��j���������   ˜wu   $�8|�g�'?�I�D��4�dj���HP�F�s���Y�*6��  �bw��z����Hg��)���l\lIܞ�����   ˛�  �������0����E�777�&�����+���g.Ǖ��x`�ڨ��  �b313�������*������dQ�����  �;  @J��db�O��H�RQZ[[s�����bwuh4~������k���   (����>�T&��***bŊ��'�`����  �;  @�J&�?��s��K/���l����\�>99��T:�=~.6t��}�DU�#  �p%S��J��l��(//��+WFYY٢>W�  P���  �������gff�tttDLOO$�����u+c�   (4g��Ǒ=���d��=�ۓ�}1%����   �;  @�����E�/��bQD�%%%��ٙ��g�$���%��?8s9��ƿ�zK�UU  �rwcj&>8{9�G��J29}ŊQQQ���M�ݻ7   (Lw  �"PWW?��s����d��r���+z{{#�J$�����|<��veܾ�#�a  ��&;7'��Ǘ{#��X*���$n���Z���  
��  �HTWW�&����gLMME��"r���t:�H�3��sW����x�ֵ�T[   ����T����/���ߒ����;w޴�V�^�?�x   P��   E$�tL&����Kq�ƍ(t�����g2��/���+GN��kW���]��  y-��~�Ӿ8z�?7��R����3jkk��6l��~8   (|w  �"SYY���_~���BWQQ������E�|I&��#���k�����V���   ����x|p�r�M��������_��%A�����w_   P�   E���4�}��x��Ws��]�1�=�������x�/'��]�u+��4w   �?{����8~u �Lm'OtttDcc�=/�۷o�۶m   ���  �H%�������q�ҥ(tI����-r�+e���蕾�28ݶ.��  `������^���T@�H&�/fܞ�������[  ��"p  (r{����{/Μ9S�ᾘ����/r�+�NN�k��[��������4   �l:��g��䓶��hjjZ��%��y�X�n]   P|�   Ď;���>��|�^UU%r�k%�N�^������n�խ�w�  ������=1�J����hnn^��%[�x��&>   ���  ��{�'����w����>3>=o=kښ�lZuU�  0�Ʀf��D�ȍ�|���---������x��'���=   (^w   ��֭[s����[�{GGG���͹28��c�uMWl[�e��  p�2�l��?�^鏬���dj�b�����hhh   ���  �/ٴiS.�>|�p�O7������N�;�R��]���G��n]�u  �]]�MmO6GA>jjj����E{^ru������   �  �֬Y�����_�"��t�$rO&�_�vM�ο4<1�}x26t��}VGU��  ����MŇ�z�|�`@�J�����E{^�<x0*++   na  �J]]]��3��O��H�RQȒ�T�;�F�\��nY��숒��   �g����<�{=�*������E���СCQZZ   ��;   �TKKK<��s���/���L�$rO.p�_�.r��I�������q��k���:   ����T|p��gN�$6O ,����ػw��  � p  �k%��?����_���¾�������I��T��x�r�xܶ�#��[�e.� ���t&>���z}���W__������+V��ݻ   ���  ����:����=7�}ll,
Yr����md�sq��Z\�{7����-  ��Cq��՘N��]r��յh�۸qc<��C   ���  �o����#����(d��n2]opp0�ۘ���_��kچ㾍k���"  ��1:9�?{%����Ŏ۷n���sO   ���  ������s�=o��v�;w.
YCCC��M&�[%Ϸuep$z��b˪θsMw���  P�f��8��@��:Y�!Y&3n/))���/n���   �E�  �����Guuu;v,
Y]]]�O�;�E&���W����Pl_�26t�  PX����ǑWc:�X.��wvv.ʳ��=�X�^�:   ���  �<������|�AA��"wn���l����8�?�mX-u5  ,��������T�r��������سgO���   |Sw   ���[���Y���[��f�P%�{�J�ڵk"w������_N���ָg����p,  �Q�!�/�������f1��d�߁���6   ��p�
  �MY�vm<��3���<R�T��26Y�=00 r�;K~w����hܱ�3�X��%%  �L6'{��'W�"�)�yS�������mQ����IܞLp  �o˻I   nZkkk<��s��$����P��Ԉܙ3�t��bO��Ms_��  @��:4<%Ƨg��Ōۓ��'�|2JKK   ��;   󢾾>����_��}tt4
U�wuu�"�l��>n���t�}�\�nm��6����   ����t�����X�3n߰aC<��#   7C�  ������Mr?|�p|��Q����s�{�ȝy���h.�ټ�=��neT��  �tfә��ro��n��Z�u���eQ��}���뮻   n��  �y���~ꩧ�wމ���lPUU%rg^e?��r��Z\�>�ׯ���  ,��������K�1�J,g��'gA?�p�_�>   `>�  X;w��8r�H�$r���>�;�fr6�=u1N^�{֯���   ^�ȍ��121�ܵ����eZ�?���bŊ   ��"p  `�|��ߏ������]�xeee.rO&�g2���28>�?9+��ލk���:  ��7�������t<�,V�^QQO?���<  ��"p  `A�z뭹����_�t�0׻�'��E�̷d��GN�Ʈ��{튨��  ��%ۓ>��g�cnn.`�+))�����9�B�������D   `�	�  XpI�}�С���~�T*
Q2�L��B���ř��q��Pܾ�3��銊��   ���t&�}�'{"��S3nokk�}��Eiii   �B�  �(ZZZ�?�a����199�(��W�X����ҙl����㮵+bSW[.b   ��䃣�>���zc&U��(N��®���T��~Κ5kb�Ν   I�  ����������w����M:/D���I�I�>;;�&gS����q�Ӂ������%  �����8r�'Ƨg
I2E=9�H�\ڝw�۷o   Xhw   Ur������݉w�՝&���}߽bv�I�b�	�@�!��Lz�O�+g:�L���B;�m�b�1��}�U�kL�ɮ*=�9�|�RUI:ǖ�[�{����q���(GUUU_���'�<S�q䃳�?8��]͍  ����8������������u�{9O<�D�ٳ'   �fp  ��x��'���#�y�X[[�rs�Amhh(���6���t�z�����mۣ��6  `+��_�?}v!7�C9J;�m۶-jjj6��������  ��E�  �[f߾}������Z���D����������Ym�l�φ����Dܻ�7����jo�  ���/-�{��K�Q(��Ԑ������@�o����x��7�!   ��UN   n��6���������oY6���{OOOnt����l���x������Hܳ�'��苚�  �r�����σO_��B!�\����p{U����҂��>��   7��;   �\KKK����9����QWWWnV��WW������H������*�  ���j!N_΋<�VV�YCCC���oz���{�G}4   �Vp  �(�������x�7�̙3Q����r����X�Ͳ��'>��b(��������  P�R���K�yQ���9/����������+l��{,��   �[I�  ����3�Dwww=z4��֢ܴ���0���hY�|��/��^�v�}]��  ����<�K��޹��_Z�
��w===�nO����?�C�:   p�	�  Pt���������B�妹�9�܇���ܹ�f���ˍ��v�Ǟ��Mo  �U(�ŧ#��޹�1���U��GR�f������?�G466   w   ���ݻ�����������Qn�E㴵���PY��)~�s��ӟ������bwOG  @�I��?��?}v!���onߥ��=���6�k����O~��  @�p  �h����/~�r����r������ҥK���p+�����F�C�]���5  �|16�����[MjmO�����o�'�|2   ���  P�jjj���������ܹs�������~r_YY	�UF�g��?������mۢ��9  �V�81'>�"�f��z***���7��7oN���������   (F�   ��M�s�=G����{��B�)�?00�C�KKK����L��އ���-��=�M  7Å�x��`^|	[Qz����/7�kTUUŏ~���>   +w   JFj���#G�D�P�r�.0���CCC1?���[�<zۚcߎ����  �����>���s[Uuuu�᭮�nӾFCCC�����d!3   �M�  ��r�wFwww��W�����('W�!�����b049oL~��ͱo��;  #��ua|:�=w!�f,�ek���͋�S�}�������   �N�  ��������J���188�$��S�?]Ԟ��(CS3���Ggsc����{:  �U
�>:��bL͗עe��U=5�of�����Gy$   �T�  P�҅ߗ^z)�~��x����ܤ
��6� �b163G>8���;�bOOG^�  ߥPX�OG����y���b ��͹Y}��T齓ÇǮ]�   J��;   %��������7ߌ���('�Bw�=<<,�Nљ���ߟ�4�����z:�R� �o(��e>��Z?o�l�������6Kj���O~��[   �R#�  @�۳gOtuuſ�˿���|������*� ?�arn!����B����%� @�ri4���`�--pYjkO�a���fI���?�|^4   �H�  �����/��r���188央�.�ҥK��,Bq�YX�?|t.����w�DU��; �V��Z��/�Ʃ���R�=��7�U}߾}���   �2w   �Fj&{饗��ߎ��?�Iuu�W!���ŀb5��<s>����;�����*  (o��+q����ɷ���Z������7��>;w�   (u�   ����ƿ��o�P(D�H��s���\@1Km�)��qGog�7��  �%�������xp4V�h����&/ZO�͐B�/���6�  ��$�  @YڳgOtuuſ�˿���|��+ۙ������T@�[^Y�.ǇG���ط�/�7�� ��glf.>X?��th,
kk�muuu9�^�I;[������(   ʅ�;   e���5^~��x��Wcpp0�IgggTWW�;��z:si4�����o{_l�l  J�ŉ�8}a8ΏM�����o���<�@<��C   �F�  ���."���K�?�!���X+�f��Op###e�sQ�R(*���Ƹw{o���Ȼ  P��b�O�����brn!�����-���7��{���;w   �#w   ���{,�������B�墩�)7����j@)���ߟ�4���bܻ�'���Mj6 ��-��1>�4��_���� ���x���+�7C}}}^ȟ�   �r%�  ���gϞ���_��W��P>��uuu�m۶�t�R,--���������_���==QW�m+ �[e~i9>�.����J W'�"��766n������s�=��   �3W
  �R����W^��^{-���X[[�r��'���ᘛ�(E��+������ξ��o{o4��  7���|���p|:<�By̕�f����������
�o߾x衇   �w   ���t��/ĉ'����erO�{{{cbb"(U+�����p��8�m�q������  l�4������_��&�v���9ܞ�o����x��gs3<   l�   lY>�`�ܹ3~��_���b���R�.�����Mx��)���81�GkC}�=�w�wGuUe  pc�WV㓡����P�,,p}Z[[���;/:�hy��f��  @1p  `KK���_ƫ�����Q.������CCC���P���g�ǻ�.����ս�^� �Z��/��ǗF��9��K����My�{�����   �"w   �����x饗����q�ĉ�i=��������t�R,//���4����8}q$�ۚs�}{gk  ���gpr&N��G���Ƥ�z{{���i�_���*�z�رcG   �V%�   _z衇r ���^+�@xuuu�����c~~>�\���ŉ�<Z����;��* �����O���C1����K�������|����Ə�㨯�   ���  �/�0��/�����s(��f���������r35�<s>�=w1���̭���� �U��/��ǗFce���H��nO-����<    w   �+����ӟ�4�z��������Aggg����{��L�RC����ő�ok�A�흭 ��s��ə8�~>t~l2��������QQQ�������]�v   p��;   |�Ԝ�.0���뱲�堥�%o����M����81�G[c}�=�{z:���[a @��_Z�O.��G��1����koo�����4G��O~���  ���   |�;v�����կ~���т���144����lrn!�~�y;s>vv��]��1��  ��J[�G�#���P�Cl����������m�����SO   ���  ��H�������~;���(5559�>22sss宰����Z�o���aw�� @)Im�g��r[���b �'͛������vC_7��ӎqw�qG    �+x   p�<�/n��曱���.]T���������[Eju?��x���Z�����n����<_���������)��   PN�  ��ٳ'oO��_�*fff�����f���^(�
�� @1���F{{{tuum���޽;:��   ���:   �F�i���E����q�ԩܨX�R����@���r�V�� (����I��}�����>��q��w   pu�  �:<x0v��o��FY��S�{
��&������蛭�w��f���  �,sK��ɥ��xp4f����|���?jkk7�uSX��^����    ���;   ܀�;w��/�����cxx8J]j���������R���O>�cg�Ƕ��t��վ���"  nTZXwq|:>���c��K;�������F����{�'7�   �N�   nPjx��OǏ�'N�ZS����ϕB��B!`+Ka��c�y�&���qWwt�4 �����3C�qvh,WV�u��ۣ��kC_3��?���y�4   ���  �y衇���o�W_}5����544��CCC���@���j|48�G[c}nu���;�k�� |��ť8;<�\���� n�+��555m�린�/����   p#̬  `���_����o�ٳgK��=5ϥ����HY��a#M�-ĉO/ğ>��m�q{_W��n����  X-��c�qfh,���r��	�A������]�6JEEE8p ���    n��;   l����3��'�|G�����(eW��&''c||<��Ka���y��:��o�����  ��t^0<=g������X.� ����������܍�Z����hii	   `c�  �&��;r��������h������p7<<�B!���������X��t�}]�T�q� @�]\�O�����ј^X���׺��6�5w��O=�T    K�   6Qj����~G����{/7:������O!���� ����B����x��`����ή����� ����872��ڇ�f(NWv%KM����*:�v�
   `㹚   7����s�[js_\,�Fǚ��r���� �[Z�ra|*�ʊ��������TU P:�n-�Ǧr����T
����]]]]����y�F���^x!�p   lw   �IRc�/��x������Q�***���),���B!�������&󨪬���)쾫�=��? ��������L|24�G'��s�����DOOO��n��:�����?�A    �K�   n��5zjz;u�T��(�`xsss����R W/�宄ݏ~R;����z��ܘ p}R����t|6:�F�ce����a+I��lO�ՍR__�>�l^�   l>w   ����;w�W_}5�����������ctt4fgg�vK+�q��h���v��Ѳa�� �w[[[����8;4�����@i�������|�(�v�Ç��<   ps�  �-��K���G����{/jJՕ�����t/�n���7��Ʈ��������@	 \v%�~nd">��� JS�cwwwoX���:~���m��   ��%�   �������;�����_�7��-�SS���P�����[\�.��R_�����jn�� ש��C�3qnt"ΏN���r �+�wuuE[[ۆ�fooo��G?��&x   ��	�  @����m����⣏>*�� ضm[nr/��>���x���<�j�c{g[���-Q)� �i����q~l2>���e���&���7,����}�Ѹ��   �u�  �H���{�'~�����B�������D]]]����t`����J��4�G
����Ďζ���5UU D�����L|6:��L���j 壩�)7����FHϟ��<�   n-w   (2}}}��+�ěo�gϞ-�pxkkk�ʊ�L�)����xU��1���])���5��`kI���s#qa�XX���MEEEtuuE[[ۆ�^
�?��ñw��    ��+\   P���g�y&>�����oKKKQ�R�}۶m9�>??��Y-���d�|�y��6Ů������u� �hvq)>��/�����v�v(_���yQx}}���^sssnmOG   �x�  @۹sgnsO!��>�,JU
����DLNN�t+=����lhr&�cg�����꾳�-Z6& ����\^Е���Q�V������y~y�R�<>�`    �G�   �\j�{��⣏>������������=r�{)�PjR�}xj6��g�����ho]-���-��n<$ �i�P��RK�����[Z`kHa����hkkې�KA������   @qp  �q�]w��ݻ��^�K�.�lz]]]l۶-FGGcvv6��ofa)>ɣ��2z[�r�}Ww{4�� ���Ÿ81_�MŅ�(������ڼX:ި������'�   ��	�  @	I�_z�8y�d���g
�(EiK������>66V�?�����)<��Ϝ�������;�ڣ��9*+* n���ZM����ߤ�G'cj~!��+5��yc������Ǐ~�����   ��	�  @	ڷo_n�����܄^����s�`xx8��R[��󨮪��������;Z�Q�; lay%�������ӱ����VUU�����ظ!��cǎx���Bk   �4�  @�J���������ĉ�������:bbb"�x��r�0�Ԝ��ܘ��;:��o7lH�& [K���ӳ���ߖ/ƧbrNK;���._)ܞ�7*���SO��&   PZ�  ��=��Cq��w�o~�nsooo�m�###���@qI�hF�g�x����������-1��]-Ӱ	@�I��\���cp},�hi�.-�Ls����y��۷km  �&�   e���9�����{q�رX]-��P
��v�ԟ���x�v�+a�q!jk���9�[b[Gk4�� [���rO����}n�c�oSSS�[��|�F��l���	   �t	�  @�������_���RTUU�����166�[������4���{-Q[�H�r���#�s�����T�����hii����iZ��;�����   e�U%   (3��^�ӧO��o�+++Q�R�!�,��ñ��@i�YX��������ln�����oo����\��ҴZ(���l�M������_,J��;�;R=�Ӽ�F566Ə~�����   �<�  @���{bϞ=��o�_|Q�M�i��������� JS��3:=�������2��Zrؽ��):���X
��L����l\����X-�޹%P��ꢯ�/��nD
��ݻ7~��    ʋ�;   �����x���O?�#G��dzn~���m�###Q((m+��8?6�G��͍����U轪�2 �5���ٹ�����}6��܈4�kooߐ���������i�   ���;   l��v[�ڵ+�|��8{�lI���m�o����177@�HA��L#5��6����ii�z�h��� `s,,��]6��f���ͭ� %�������7"��?��Cq���   P��  `�HA�g�y&���_����(5UUU9133ccc�ܡL�Pe
Z�����|_s}]�v����[Mu����_Z���hj&��g��[�����]]]yNz��������   �O�   �����x�W�w��]|��Q��v�)�022R�A}���,,�G�i��[��r�=�����(�𷤝{&��
�M����R l�������ɻq݈������;�3   ��A�   ��Ԝw�СػwonsO��&�%RXzz:�����uL/,��ɥ��qMUUt47DgSC��6G_{K��x��zR;���|��\nfO��+p3�E����9�~#�^�=�\��   [�w   `K��_��q���x��J2$����U����b [�����v������|_cmMt67FWKc��6�������r��Z��ٹd��_�83�ف['�Sk{SS��N
�?���gϞ    �w    ���w�uW��7�����(5555100��������$sK�176��.�^����ֆ��ji�M�)������P�
��7��1:���=5�;��Ecccn\����ݻw��*-L  �-K�   �����������s���;�������-r��Ғ�R��Rtrn!�3_�WSU����Ҕ�񽥾. n���jza1�G�fcd�r�}�P�b���]]]���zC���O=�Tn�   �6w   �k����~�ȑ8{�lɵ�����6���>55ZM�ﲼ��&g�"��[뢭�᫦�|��"
l�o6��������Uav���Pz
�WW_�e����������    p   �J
'<��3188o��F���E)��������Hm����p�R�}tz.�+M��W�j���>޻��r�{CmM \��啘�_ȿ_R�=ڧ�-�JN�suvv��nDj~��g���>    �p   �U���+q�ĉ�ӟ����QJ���b۶m1>>����WjX�YX�����W�7��D[c}]-M����u9�l])�>���s��}�򢙙��_��(})����55׿�/�՞x�رcG    |��;   �w=���q�}��믿�[�Kɕf�������� �(sK�y\��^�h8�W]Um���P�U�=}�\_������L�/���|nb���|�\?����e#Z��k�~�����Geee    �-�   �UI-}/��R|��gq�ȑX\\�R��۷o��������Ͳ�Z����<�ReeE4��F{c}�75\�7����������A������[�;:��ف�`#Z�[[[��g�����    �.�   �5ٽ{w�򗿌w�y'N�:kk��Jm����###��� 7K����i���B��ښ��ޯ��;֏5UU�<K++1=��C�s1�����t��QR�z�C�Hk{uuu8p ��    ��   �5K!��ƾ}����_����(%uuu�m۶�䞆�p��--�qqb�k���TGs}�������߷/�k���3Ky��t^tr���# ����===9�~�v��O?�t�C   \-w   ລ�����ş����農��"�����H��E�6��� n��s�����c�u�_��S����1��������斖�
�� ����'L�-���j ��R���+Z[[��5�<멧��y   �k%�   ܰ��/o7�ȑ8{�lI5�������@nr���m�@�(�����2������ʊh������M��9��T[�o7��)U�)����w=�M����ا�����\�������������~<�@    \/w   `C� �3�<�������6fgg�����}�澰� �,5X��oߦ��:��Gcm�W�)������6��fJ7ҮWB�)����q
�ϯ�N��P� ;�ƪ���m�)�~�����駟΋�   n��;   ��R���_���?�=+++Q*jjj��?==���Q(�\�q�siQ��_}���"R �.�kr���.ꫫr8>�S@�^<W!��/,_����������]LA���ʞ���jii����r�i���Ç���7    6��;   �)�����{�ȑ#q��ْjZM������>?? [Q���ڳ�����������h���������>௄��ǵ�I�Uė�Z�_Z��F�W
�ǥ���K���_������ (*i�ojmOs��������   ��$�   l����x�gr#�o����Q*��������9���ۭR��pU!����Z�k�*s�&�禀|uUU>��k�/�_[U���iԬm����K+��c%ԗV�o�p�j�?���r`==���Ws��PB�� �������^YYy��M�v������   �=�   ��K��?��O�̙3��[o���B������������v�ƤP�\j����W�O����c��J𽺲2��t_���]ݗ��5_�_��c��</=��2��ؤ0���JnL_Y-��k��j��K���5O�IǕ��Ǥ�.�ϥ�/����W�})��b���SWW�[���Z���in�1���   �fp   n��o�=�'Nğ���X]]�RPUU�C )̑�ܗ��~C1 �#��WV�n��K�o�������7�V��W]��-���_o:_K��o�˯�`3���J����A�kU[[��n�-    6��;   p�=���q�}�śo��ϟ�R��ܷm����y��" �mq��C� �#�J������~i8���8p�@�   p3�   �D
����122���Q
R�a{{{�������|   ����loll���yO���駟�s7   ��I�   ��R�����ԩSq���X^^�R��"}}}177���  p��pzkkktvv^W�z
�>|8z{{   �Vp   ��޽{��{����w��G���Z���H�����155   �JCCC^D\[[{�ϭ���Gy$��    ���  ����:>�`���1<<� }ߩ���9FFFbii)   n����<'I���*5��ڵ+�Ů��   `�	�   E���%~�ӟ�g�}����cnn.JAjIܶm[LOO���Xɴ�  �+͟���r��Z�����Ç���)    ���;   P�v�ޝ�ɓ'�رc���� Ls�}vv6   6Z]]]twwG}}�5?7�>��OD___    w   ���۷/��ݛC���_��B!�]jOLm�)�>::Z2�|  ��UVVF[[[tttDEE�5=7�:�����w�    �J�   (	)ı�����������Ν����(v�Mq۶m199�G)|�  @qJ��]]]Q]}m�y��{�7y�    (v�   @II���=�\LOO���K��>4�Z���se||<fgg  �j���Ewww^@{�v���ʋ�   J��;   P�ZZZ⥗^��/Ƒ#Gr�إ�Ş����������R   |�Լ���mmm������8|�p466   @)p   J���@���?��?�8���?���B�Ժ�m۶����A�B�   W�]�������r���=��S9   P��  ��p�w�q������+++Q욛�s����d   ����������������k׮    (e�   @Yٷo_�{���[o�G}kkkQ�*++s�b
��6����   ������؞دEMMM<��Cy   P�  ����!�����Ĺs�>�B)}}}177����@  ܸ�赭�-/|�������ٳ'��|   �\�   e���>�{��#G���x�kll������������  �/����Օ�^��ߵkW����   @�p   �^www��?�c�����b�+�����ԔC����  �����<OI�r�Eoooޭ*�    ʕ�;   �e�0��~������㭷��-�Ŭ��*zzzr�=�򗖖  (]�?5����\���\��'�̍�    �N�   �rv��?�����O?�w�y����q۶m��}||<VVV  (���y�jGGG�}5��N���9؞�   �U�   [�m�ݖ��ӧ��ѣ���Ŭ��)s bb"
�B   �-��wvvFu��_�M��'�x"?   `�p   ��{�'��'O����cii)�UjqL͏���199SSS���  @qI�S�����������Ӣ��<   `�p   �Ҿ}��HA�cǎ���r������� ���cvv6  �[���.7�����J�ݿ�a
   `�p   ��r߻wo������j�������ɭ�)辰�  �͗�������ժ���Ğ={   ���   ��Ԑ�~�����������������n� �r��)����W�����x����{�    �N�   �;\	����[o��q
�(V�}����������� @�kii���Ψ���������~���c    ��;   �U����C�Ł�w��]�;w����)h���SSS9辶�  ��hjj���X��q<�@    |7w   �kP__�>�l,//��o�]ԍ���֖�����133  ��K󁮮���������������   ��p   ���15�?��cq�ر8}�t���F1�������vOm�  \�T������W����_�   �:�   ܀\9x�`�߿?�=~�a���D1J��������sss  |�t���y�������#�ĝw�    \w   �P]]���>�hnt?u�T��S(���7s�}~~>  �������ۣ�������?�p�q�   ��p   �@�����=�[�}��8y�d,--E1�������t����  ��,�ӎG)�^QQ�M�ohhȍ��~{    �1�   6A
�?���y����'�:���ߟ��SнX�O  �,��=5��p��ۛ�����;v    K�   `��۷/�ӧOǱc�r�����4���bbbB� �����)ԞF����f�G}4�o�    lw   ���{��#�S����l����<����WVV  �IjaO���������---q���    6��;   �M��A��Ǐ���b����U�=5�� P�RX=���`{UU��}lWWW<������    ��    �ȕ����~��crr2�M
�477����t�WWW  Jɵ�SS{jlO��    �\�    ��m�ݖ���x���;q�X[[�br%�>� (W�c��ڢ���/�VVVƮ]�������    ��p   (��/���\��f�B���/�� (V���^SSw�qG8p ��   ���   �Lccc<��ӱ��ǎ�?���B�W��i\	�///  �J)�~%�����������   ��!�   P�jkk�����裏ƩS���ɓ9L^lR�{�y>�S0  n�fokk�㻂�i�fKKK�߿?v��    w   �"�:������ٳ��}rr2�Mj�LC� �����*7�_M����3~���#    �K�   ���ٳ'�������������(&W�����9辸�  ��R��Jc{
�������lO�   P��   JP����?cjj*�y�8�|
�(&y,,,�{: �����Ρ����]����;�3y�|   ����   ���=�=�\����ٳgcuu5�I}}}�� p�jjj���=����3؞X����o߾    �4	�   ��"?|�p<��q�ԩ<�����\	�/--���d���  |����������;���?�p�ر#    (m�    e���2�U�q���8~�x\�t)��֢X���FOOO!�~�B!  �����hkkˍ��&��n߾=8�w�    �w   �2500/��b���űc��̙3���Ţ��:��Spiff&�����  [SEEE455E{{{^�m�����x衇r�   ��"�   P�R��O>?���ԩSq��ɘ���b�BI����u3}_)込�  l�|0����i�I�#S�}�Ν   @�p   �"Rph߾}y\�x1�?�.]����(�����9��:��� @y����S��ۚ���۷o��<    �O�   `�_|1ɏ;gΜ����(�u>�p���*��y  nLmmm����i��=���΍��~   �<	�   la)D��O���8u�T�<y����uuu���9�>==]4��  \����hoo���&���P�Ν;   ��I�   �܊�o߾<.^�Ǐ�K�.M����::;;s�畠{�P  �[jhojj��������s��۷ǁ���%    ���   �����x��cnn.�;gϞ����(UUU��3�R�|
�/--  �%����zkkk^����F�;�37���;    $� �����X]]��}��t��jjj�   nLccc<��y�9s&�}���b��@����H�tO�w  n����lO#��}S
�www�������'    ����TW�&i����Z Ә����15B.,,��z�/��7"rR>]TI�ߦ�{���O����k��I�Bi�0��,  [��ߞG1���s��������<�(
 �͑�������jz��o��   �Ւ�ຬ�����dno�����������P����-�>S�&I!��q�L
���LGGGy;�� `�(�V������=���r�{1�I  �Y:�J�P�VY��v    ���; �*5������p}uL#��WVV��]i���Ǥ�tq&����<��N�  (W���D�B�4��*��  l���N
���ν�I[;    7B��dO��.�ŋ�1���b�Q�����Mi;ށ��ضm[>^�  �E1����UZ������N)��@  \���ޝ@g]������$d���"��	�E�E�}��V��ڱ�e��z�̙qڞZ���.ETv
HQED�N�	KH H��^�FDH����ޯs�yB�&3��w���ύ��wm��y.��     �-� �TVV���ڵk����ݰ`�W_}%x߉'\��FU�d��֭[�ѪU+5mڔ6#   �@mu���t7,%%%�6w�3  �8{���v�ׯ�ݭE��  ��a�V�gE���io[�r	gΜ9��<�_�=�۳{UVb���_��3tt�  �7� �lc-�(��u^^�kg����l��}�v7<l�زeK�i����  �`U��ݞ{7l���JHHp��ɓ.�na��@   ���Â���n�PUY8�
<z�꥔�   �O	Gii��=�n��[���x^-�^Wl}��U_=�JDl�`���� �[�@�ӹ۶ms�O��އ�`�sC�6�ݭ)33�I!   �N�v�ܰ֠��׻g^���7;dڸqcw�>�<��  �3�[���%���h�;u��m�   ��ٍ�TQQ�>|vX����׆'`_\\\�����d`mX����4�k!x  ���; 1�[;{nn������$5c'�?��37�m*edd���m"�kTT�   �``ϳ�{�v�6w֭[��{��kt���Y��!;xj�I6hu  ���y������۶�تU+��?Pll�    ȕf�����ڰP��9r$,���ކeW������.��ym֬��6m�� ���; ;�kA�/��҅����#���$=-�,P���]��ݳ���Fӹ�   ��Q�F>|�{�n�ڸq���{�c�.�,D�;  ejk�߳�^�z�I�&   �WZp�����s�v������q׮]n�+99مݛ7o�^[�hᆭ� �w p�w�>h�p����0o޼ٍY�f�)�gee�K�..�   ��mۺa����tZ�ܟhu  ��Bm����;�5F{   ��[��ؖ��f÷��ކec<lNbn�{V�g���  �>� `<-�6lp��C�	�.�Y��c'��u��6�lc�M)   ���(���ۍ��b7/�$���  ��kk�P�=�dff���/Wll�   �pa�j���矽I�u��a<������ۼ�}����֭[��L���  �� ��#,���矻ӨL��-��ނ\�R׮]]����-<   ���4:Խm!w��M��  ��kk��Gzz�z��ƍ   u���w�^mٲE[�n�Ν;]����ѣ���O�0�}�vw�_v�e�5..N ��F� ��B�_|�{����J�d��V�X�M�սW�^43   �y�����6�({������ǏwAw�*  ����			.�~nɅ=�dee��  �Pf�vkf��D۶ms�x=v���������e˖.�ޡC�j7Z �w �Cv�w͚5.�n��i�����0m�&Wvv�ٰ��t   �@�ZFm��jݺuڳg�_o����٨��PYY����   u���4h��~��Ђ�ڵs�:��   �������{vhOv�a׮]n,^��͗����Z���`0  �� |�&L"�P�ƍ݃4H,�~�z7<�����S��ݙ�   `%''k�С�m۸������'O����d��IIInX���ݭٝ��  �W�fF�a;;xW������֭��   ������Kw룽8���Z��kx��?�[`׮]���. @�!� >`M}j_�z���܇`Q��ݚ�z�쩾}��}���T3   �5jt6�~���<�o�>���,Tf#55�|�Vw�  \*+��@{bb�ق
[���7o���vc�   �Pd!v������@M����ؘ>}�[_���6hw���wc �"P�Z�J+V�p� �Y������HIIQ�>}4x�`���	   TM�4�����ۻw�v�M���Wee�_>���Q��f��6_d�  Ԅ��[������ξ�B�-Z�p�1�   �v�ڥu����>s�����%K��a�Ν;�2�.]�(::Z  � � �Ȯ���v��ٳG@(:|����kѢE�ԩ�����/����   hn�[��5�ە��`��֦j�Z�,�ns�ӧO  �|,�nm�6<7,�3Ezz����>    Y���O?�'�|���`�qڿ9v����z�r󯪇� �G* j)??�5[[c��S���X�;�l�aÆ�Y�f   �'�nϴ[�n��͛]3����111nXӪ�m�8qB   �hM�j���t��ڻv��Z   BV^^�>��cl?r� �,���ذ9Yvv�~���2@[� �w ����rwJ�>��a�N.�!�?�PYYY4h���y6�   �@T�^=u���O���/�t��#�nM��VV�|�9��;  �ǚ=�����;סC��   ����b�Y�F}�M�Xg��f�~���fw� ��� P���ג%K�z�jr���溑���������L   ��j�����r��URR◰�}>�`[ee�������ɓ  ��B���n��ƺ�YyD�F�\��]�v   Bѱc�\S�e0�������6��V�+��Bmڴ �{��l۶M,���k�`b�Ľ�3g���>\-[�   袣��3�O���͛UTT������Шk�4�v  ���x;�V5�nA���t�o�^m۶   �l�mӦM����׻5/ �ٚ�e��hڴ�������6 ��p�sXkߪU�\c{AA� Ԝ-F�ב���,6L]�vUDD�   �@W�������e�wE�?6�,�f"6��ۦ�5�[S  |�lѠAl�W[#���7V�ΝբE   ����>��C��~��Q�j����9s�f͚�.]�h���֭�� j��; �����裏\c;�*�{��k�2d����JEEE	   ��`M��6�ݻw��[ۘ�G���ᒒ�ܰ���naw�  ,UC�qqq.�n7�4o�\ݻwWJJ�   �Pe�7ntł�����6lp��q�����+--M ��#� 암����/^�'N�oj���?��_}��ns   &n{���/��_��OZH�Frr��[�����J ��g�v[���n��Z�r����   eV&h�|��:t萀pg_V��p�BeeeiРA�ѣ�� P��-k۳���L�P��P��ٳ�t�R:TW]u�{   JvK�cϹv���w��u�J�Fjj��fw��:uJ  �w<M�e����H%&&�P�]I+    �mݺյ���g�����zqnn�M�4q9�+��­� Ώ�;��STT��}�+��,lcA�E�i�����԰aC   �ȞemC�Fii�>��s�޽[ǎ��ϥj�����ݭ�  \����0{�P{JJ�ڵk��h�  @8�u��������v��! �c��S�L�;Ｃ����ꫯVZZ�  �F�@� �&��i~��$�  �P���p6�n�Ok�ڶm�����Q�x�|m�6O�8���
  ��~�Z�݆��GEE�q��j߾�233	�   lX��|�e˖�[�Nyy��J����_��vp �5� B^aa���}}��'u~E<��t�븮��w�3   �,�ֱcG7����]�}�޽�U�.Y0/11��[��vg� �wY���Y�ݮ��ז-[�K�.��   @89t萻���s�)�[�]�v�p���kյkWEDD �w !ˮ�����ŋ]K��`�!����?��O:TÇw�X   @(hڴ�櫯�Җ-[�ζAXYYYg���-�g���r����r�  ��:Tզ���T0���hi  @X�R��K���[��om߾]/���Z�h�J{����H@8"� �؆��\t]_��{�ky����j;�6�5N   �"::�5��0�����w=m]��[�ݞd�>�}lO�;�� �Pg����8�s�B�v��y�����v�v    \���kΜ9ڰa��u�n ����{������O^@����aavkk�?�ۄ�6��3gj���=z�z���U\   IU��-dna���<>|�N���a,�naw�9 
,`av�/��m�ֵ��4    ��ٳGs���ڵk	�~V\\�I�&��I+���+% �=�P����EEE�<�q��)33S��r�ڷo/    T��ƺÝ6N�>�;vh۶m����������6t���v�܆�+++ @0�\����Ҟ����eee�q��   @�dV�2}�t-Z���;��A�@P۹s��~�mm߾] 5X���U�n�t�m��Q�F   BY�z��O�!OkR���]m>v�Y]�p���6--��=�w�� ��iٍ$�s�j�Ϯ֭[��   �Â����6l�  ��j�}Ĉ�߿�[?�PD�@P��3f��� -����jذa����#    Xm�.]�0��a�wی<r�k|��a-��1������  @UU[����բEu����   ��Y�b޼y�裏X����	���[�օ뮻Nt% J�*Z�l�;=|��Io�T9�|�Z�J7�t����ˤ   a'%%E�{�v��߿_[�nUAA�JKK��Jik	��`BB���5�{��� ��ii��Av�_��͕��ō   �;v̵?/^��e0 /;�2q�D-Y��5����K *���<m�4	 ���ʜ�}�ᇺ���ղeK   �iӦnk��������u��A<����5�ڰ�}r���}|� �ڲUh�a7��P�6mԶm[   �0[����\㳭� ����+���}�|����� ;� ^aa��N��/��B p!�R���k���5j���   -��	����m۔����}���ׁ��aDSYY���w��  ��n�S�3$99�m�[����.s?_    \����^�Z3g��ѣG tmڴ�e&z��1c�(--M ��X��m���}�]�� T��C.]�T�~�������O    �f!�.]��a�6$;(ZPP��>u��?���H��ǻa,��	�۰gz @����9hoѢ�Z�j�v��)::Z    j&77W3f�О={ <ء�K|���:t����z�. ���;��dmr�&MrW� @m���(''G�|���NN&   �a��޽{������6=:��V�~}%&&�a쐻���^}�0 �/�9РA%%%�u��n�iӆ@;   p	
5m�4mܸQ ��W_}��F��>}����  XpP�������]+V�`�Wآ���iĈ��꫹�   ��sޭM=//O���:x�JKK}>_��^t��o!wϰM�  �EEE��������왙���    ^�	�ڨ��� >����^Ӓ%Kt�w�98 � �]�3q�D�` �d�vx�N&�;�m�   �8�m��c��{�����\ི�ҧ�Z}m����݆}N ��e�v�>n�v�D�ܹ��4i"    ޵a�M�:U����sٚ���g���W7�|��5 Pp�wǏ�̙3�|�r�/�ٳ�Mج��G?���   @�Y�<##��4ݱc�{�>v�***|���
]k��a�ƚ�,�~��	x�e� pa�}:::�m�7j�ȵ�ggg�aÆ   ������ɓ�y�f��X�ȪU�\	�1cԿ7��@D��_}�駚2e�� ��`a���&l����[   ��IKKs�w���ׇ�Ν;����f�s_� �'Li,`�iw��u� �;v�)..�؛5k�:�P�D   �[�����C���O ����2���Z�b���_�E͛7 � ���&N���k�
 �a߾}��_��믿^7�p�ې   p�RSSݨ���z?x�JJJ\뺯�MM			n���w���c@�������n��ܹ��6m*    uk�֭�4i�


 ��m�6������o�Q111�@A�@��k�rrrt��a�?�>}Z�g��ƍ����L���   �}~������]������� �������<�B�6,�n��w �.+�&���$�fҩS'7(	    ���P�O��իW�̙3�Ke�A,Y���&��=++K ��3�@4w�\͙3���������\7�|�$    �e��mۺ�QZZ��{��ё#Gt��q��x�6<l��v�໵�[ �EDD�����a���4]v�e�޽����    0lذ���ۺ	 x[aa��~�i���W��v�4h  �'� �]E>a��� ��,'Nԗ_~����]�   ��X��s��n��z���<�cǎ� �/DFF����6�(o�O��^9� TDEE����n�Zݺuso   <�&2c��Z�J �K��i�krss]��~ !�����g���>ۄ oZ�v�v�ܩ�����С�    ��5�7o�܍�����{�n8p�5�Y�ؽ�Z�-to��控��z?u�  �U�gdd(;;[͚5   ���駟jʔ).� u��ѣz��իW/t� �?p�36�z뭷�~�z@09|���|�I:Tcƌq�    �������j�޽ڷo�:��Ǐ{=|���X7<�e�>�O�݆� �}����vs5j���Lw+FJJ�    [ۘ4i�֬Y# �;d�}�v�s�=��� �%�Z |®�y���]� #kg\�d�����g?S�&M    0Y��cǎnxTTT���@{�����]�B����-�2ㆧ���-��	�۫/Z��/��cn���\{۶mթS'p   �v�ء	&���H �o��z��)P��n��l������zs� �%??_�?��n��v���_    ��m�ddd��a��v߽{�{���N�8���}l4����4�[�݆�[�����(w��^a���0O�-\c;   ��aks���ܹs�@@�nڴI��{�[�  _#��klSx���ڼy�  �X��7�p����.��    �X���t�Mָn�h���w�G�uW����u��Ӷl��6�-�n�w{�: �k_�� ���q��.�ޡC�o�   �l=�Zۭ� վ}���?�I7�t����*��)� �b۶mz�W�0 ��U�V�	�����Z�    �k[oڴ��*..v����B��QZZ���`����7��P�'�n!{O �^�1n��k�ݰ7�[�V�v��   a�� 'O��J�  ��:������_h�ر�> �w �l���:u��p�P�k�.������v�S�N   ��p��Ν;��t߻w��>|�l��W�[ ֚�m��j��3��qx�� ���SRRԼys�m�V�Z��f8    ��%���Z�~�  �X������]Ƚk׮ o#���l�N�X�B Nl���g�Ս7ިk���k�   �0�����;�Q��,�n�����Ǐ�u�_j����8�߫��W}���O�=>>޵��a���teff�fv�}    8�M�6)''GG� �cǎ�^���u뭷��� j��;�Z���q��iϞ=�pd���3gj����{'    ��kj>�5�:tȅ���ą����]�R������&6����s#pa���ns֚���m�7m��5�[3��>    T���g͚��r @H��e˗/�Ν;����� o ���6nܨ	&�X wve����'����q    �>��`��s����UTT����~d��'O����e���>��B��f;B�}}DEE��!��n�u��l����ccc    �`��W_}U����Pc%��?��~򓟨G��KE�@�ن��"~�w�܄۔oԨ���PPP  �8p@��_4v�X���S    PS��P�����n��eeeg��{���ǵ9��]�	�WVV������ EDD��u;�a�boذ�[�JMMu-��j    |i׮]z��ݼ B��T9n�8]s�5�����# �w �b����nM�-��g-U6�m��ܳ�mo{ެ�*>>�]�nv%�m�m޼YS�L�l���+��nЈ#�   �Uj��E���O��B!x��m6���]Y˺�m��q��JKKs�����   ���Z�J'Nt��@��u�(//O��w��@mppQ�!����+??_��gmT�a|���m���_l��:��k6Q�={���ۧ{��+_c    P]�	�;v̅�m?~܍'N� �'o�tS�P�5d۸�oYӻ��=�j;����~|�Oh݊<ֺ�Y�JIIQzz������	�   d6ǝ:u��/_. 7V��������Wff� ���� iZ��k����/��2eeei���:x�ڴi�m���&�m,�ƣM�|m�ڵ:|��~�_�w    ֘d�u�����F��G�����-o���	�_,ok�	�{T�����@`��ok��a�vd��ຕ/Xh݆�-Y�zrr�{��j    ���
Ǎ��;w
 }/|�'t�wh���� ��{mڴ�M�l���6 -�n�m۶n��t���/��m:������P �a�Uv��P�V�    ��:�����._ZZ�֒��6,_�ޮc�\7���$_��{� �������'$�ayO(�^=o��<A���m�ʚ��՚���ڍ���+    [�l����URR" w���o�����Z�j���Z�b�&N�ȕ��6-�ޭ[7l���/5jԈ�;pG�����7����:w�,    U���n4iҤ��[�����`��Z(�jS���m#�jx�s���V�Wf_���ws����x�/��<�s�����ϳn����������{�����������R���Ն5�[P    pq6�[�d�f̘!n?�y���z�ܹs�T �-_�\�v������. �b���p͞=���m@�o�^]�vUǎ]V���;�����^w�y�$    ��Y�ښ�mx���[���������m��y���sٟ;7�na�s� �6�{�/�n!����?�	�WekD>��������~�8�W�D�߳p:    ��ٜ��W�^-��ۺ��=��ږӰ���ڼ�s���y{�� ���IOO'�����|����/~�eff
 .��;���p���4j�ѣ��7v}�>g ���&Mr��#G�    ��<��6     �b�_z�%mٲE<�g�ԩ�Z�h�iӦ��zFF�Z�n��V藒����Di ���G��'�Џ�c���G �}�p�p��M����ճgO�j�J��q��pa�2:�������         EEEz���~!p4i�ą�m����k��^5k�̧a��!�|۩S���k����1b�yoD � \��g�a�����.�ޫW��^Y�l2f��^��V�X���2�w�}罢         @�۹s�^x�;vL𿤤$h�޽����2-[��?X�<�o�Z�}�ر�' |w ���'�t��Q7l�ԦMj��U(�8[}bb�JJJ��֯_�g�}V<��bcc          x�[�ε��W��X�`�Νխ[7eddl��)��O>q��_�򗊏� xp5�?��S:r��{vҰG��ׯ�kn5��N���-[����>� �4          H,^�Xo��6ae?����٭�݂����l��6�ѣG�v�ء����.?��* �C�S�w��3�<�UYu����{�V�>}ԠA�*��'�������O?�_��WJHH         ��t��iM�6M|��P��Vy����3(��� �|������ֿ�ۿ�C, @�C�|��gUVV&�NJJ��&X�pb�R�d@��ڵKO<�z�!%''         @`9y�^}�UmذA�[�Z�R߾}թS'իWO��2۷o��g�@,?���\�����af�֭z���U^^.����=z�䪦��g'���~��%          �Xy�3�<���|�nԯ__�;wV���դI����4�8˴������{]�
@�"����7��_֩S���`��\���o������         �����p��={�kذ�kk�ի�bccJ�T �WQQ�W^yEw�}�;� <p������~{ �w%''k�С�ڵkX�=�fP;�rM�=��Z�h!          �a{wO=��
߲v�>}��`����"�@͜>}Zo����!Y.@�	�' ����+''�����4h����ׯ_�N�j"""�M����+ �g-O<�|�A�i�F          �ݾl�v{��n�ZT���]� �Q�ܙ3g4m�4W�:|�p/$2��z�jn����pX���+�Ptt���w?~�]u����E          uc���.�~���7Z�j��:tP�� �5��۷O ��2o3f�бc�4z�h܁��g����_'��%6��֭�;��� |�M� xǉ'��s��7����5k&          ��{�nWDeAJx�ۇ��m�*Yi w�v,X�2pr� |��;�rss5~�x�>}Z�t������kմiS���d������O?����w|}         >����g�}Veee�wY�}ذaa{5{���Y�p����u�wr� w m߾]/���***�K����k��F�:u.�q���]v�����7�����         ��nݪ��'�=�!�����l¨���^�����t߫��իWO Bw ��ܹӝ(>y�P{����ݻ����*EGGՓ����9 �C��mroذ�          x�ƍ���/�ԩS�w$%%��+�T�=�VA�;����&���?u/ ���;B��٣�{�ŗ(33S7�pm�`��z_\\, �UXX�B���o/          �fӦM�۽�
��﯁�~}bi�wJ�X�f��Z���8H�(�$�q��=��3*++j'11Q�^{�:w�,Ԟ�8&���޽{��SO�׿��4h           ��c���⋄۽ ""Bݺu���Õ�� ����������p�֮]�7�|Scǎu߇ ��@8x�|�I����c�vkm'0z�,�y�f��ݻw���ׯ~�+���         @�؞�s�=��'O
��u�֮L�Y�f��Y���;�=+W�Tll�n��v-܁ g�O?���9"�\rr�F��v��	�a�1 ��}�v���Kz��%          ճo�>wk���ǅڳ�aÆ�gϞ4'�@ZZ��n�* ޳t�REFF�[n��A�b����DqQQ�P36��ӧ��lEGG�C���������}��ǂ         P����D���L�ۛ�֭�~����;j�L����?����뮻N Bw HUVV��_�޽{��IJJҍ7ި6m��׸qc��~�������4          �����.�~��Q�vZ�h�n�A͛7j��;�;�f�rM��\s� ?�@:s��z�-�ދ��ܹ�F����8�7bcc݉���R�y��)99YC�         ��*))�SO=���b�梢�4x�`���_���j��;�[3g�t٥+��R �w ͞=[+W���\���zwM|�&d܁�3m�4����=         8��]?��:p��Ps�Z�ҏ~�#��^b���a)// ���ɓ'���>}�@�"��O>�Ds���/33S�G�VÆ��aۼ�<��O�ք	����N-[�          ����z��UPP �LLL���^�z)""B��T�ٳG |�B�999��X��� 8p��֭[��믻¸8�ˮ���Yu+--M ꖝ�����#�(%%E         @8����+���ݻw5�����n���"�Lw���(p���z��ծ];>܁ a��_|�EUTTgW:�d���j2�?�9�g�}V�������8         �Ȋ�z�-���
��A�Q$�cd*��q��)��������t.܁ PZZ�~���Y�����k���jР���7 �طo�^}�U=��,:         ,͞=[+W���V$جY3���u�rwVh!���D܁ g'�^x�
�誫�"��gIII���r�~Խ�7jҤI���         ��O>�Ds���ǲ}����W_�������@�:x�ƍ��z��s@�`veք	�c���bbbt�7�S�N���8--M��� ����]��-D         �`�֭z���]���#G�s��B�IMMuō�O���a?rrrt���\��G�`���Ӻu�kڴ�n��V7@�����1c��٥K         ����@/���***��kѢ�n��f���u+22R���:t� ԝ5k�(==]�F���G�P�6m���/\X�4f�����Z��yny��G�$         E���.�~��q�¬�x���:t�k�X���;P��Ν��\y������X�Ǐ�*��	׀4l�0��	P܁�`�x����#��+        �Pr��)���*,,.����8;;[�/�TlٲE ��ԩSոqcu��I w ���kܸq�t1ί~��9r��w�..�@��srrt���s(         !�s��;��=��n�ͅ:�d* ������/�����wjٲ� &�@��<y�����KHH�wܡ-Z�---�imA��}��g�?����:         ���w�Ѻu��ڵ�+����e* �Oyy�^|�E=��JLL��C� ˖-ӊ+��KMM�]w��^��������Ç@`x��w����5[         zV�p�B��Y)����5d�!����_qq�^z�%��׿V��Di�@�W% 캬�ӧ痑���4h ��p���?��� 
         �8���n� kk=z�������20Ǐ �پ}�f̘��o�] w  ����W^QEE��]��ٺ馛\#8��ܷn�* ��رc7n�~���*22R         @09y�k�-//�/))Ʌ5�5k&���4�@ X�t�Z�l��
@� ����ӧ5~�xZ��G߾}u�׺k�|�RLvkȻ��         �`a����


��kժ��[;8�e*v��- �7y�d5m�T�۷��@��Y�fi˖-�w٩����Z^v�@`Z�p���u��M         @0X�`�֮]+�_vv�n��&EEE	��L8*++]I���G%&&
��p�h�֭Z�h��m��~�5��+���@�v���=��cJMM         �6m��n)�����O?��]���LX�9�B�=���ի' �E���Ǐ��^��ӧ�o���ȑ#գG!�%$$�k���;��c_�r�ᇙ�         `:tH���*��}�k��V}���w �l޼Ys��q�5 �E��I�&�	���o�Y�:uB�]�E�\[�l����u���         4�N�Ҹq�t��1���ׯ�1cƐ�R))).+SYY) ���mڴQ�.]��~��Gi͚5�7���[nQVV�Z����ݻ p�����ر�ڵk'          �L�2Eyyy·EGG��nc�/�YV�B�EEE8Μ9��^{M��\�' � �Ա��BM�6M��=��z�.\��ÕZ@೫'L���{Lqqq         ��U�\� ������Nedd��2܁�SVV�r���oU�^=�{܁:d��<yR��]�e��:���;��������'         ��B��ގoKHH��w߭&M���L��o߮��_�F���G��C�oǎ��<���C�1 x�\�R]�t�~�         �b�������˅o$''k�رJIIB�
 �͛7O;vTVV� �-�@�]����fW��=�p{���5�WTT@���.�LIII         �aΜ9.g�onMiii�Μ9�	&��SÆ��p���'�:;a����7�t�:w�,�>��NMMUaa� ���R����z��!         �.����\|�p{��|%%%z�7��_��P��u`�ԩ*..�~ȏ1B]�vM�����/�ԇ~�A�	         �+���?~�*++��Y÷��iMqqq���WYY� ��7jٲe2d� �mذA�V��v�uשgϞBx��1|f̘�nڰ         ��0e�	_������'JLLB�e*���r:tP������>t��	M�<Y�����էO!�؉r ���1슭�z�+�         �sk׮�@����$���?&�,����/ ��ԩS����#�<���H�-�M�6M��^�zi�СBx��N�6m�ʕ+տ         �bي�'
_KHH��w߭��d!�Q�]�vi�ܹ9r� �w�Grss9Y��u��Q7�p��,�n�gΜ��2}�tu��I)))         ��������L����5v�X����@p��{�.]ԦM������7� ��Z�j�[n�E����WLL��6���D �ˉ'4e����         �m�-��͛)66�5�7n�X܁�r��iw0��STT� �w�f͚��
w��{�m��~}����	w 8�_�^�֭S�=         xˁ��{�	Rdd�+lڴ�^���]����B ����z���5z�h�R������kٲe
wqqq�뮻��Y�����; 8Y�{VV���         \�3g���7�ԩS���ի�1cƨ]�vB������T
@�X�p��w���n�G�^d׏L�8ѽ�3;U|뭷*--M�Wj���ѣ�=�n�          .��ŋ�m�6A�����l!|YƆ�;\��[o��?����� �"�x�M�v�ڥp�Q�F�M�6�"���K��w��j۶�         ��***r�J����}�
�L�


4o�<��G? �"�xɡC�����+�0@ݺup.&c@��Ǔ&M�����:         ���=�7�xC'O�T��ҥ�,�L��ϟ��={�e˖�=�/�>}z�O�ڷo����J��$&&*&&F,R �mϞ=��?���C�
         ��+Vh˖-
w�[�֍7ި��܁�UYY���zK����U�^=�����jݺu
g��}��7�C��&���d�޽�f͚�^�z�aÆ         ����L���]jj�n��VկOt_#����<W8d�����Kd'��N��p�;�C���.��;���]���?��         ��>}��;�p֠A�u�]�������İ�� �����˕��, ���;p�/^����+\Y+��Q����&�b�w��:rРAjӦ�         ��ٲe�V�^�pV�^=�r�-��8�e*�����~�m�w�}p������Ds��U8�pcVV����J- t�9sFS�Lѣ�>�;         ߧ��B'Nt{L���k��@
��2yyy�֬Y�+��B]�t�KC�����u��	�+�t2D@upBK~~�V�\����         �>.ԁ�.��r���G��!S���S��?��?% �G���ݻw���Y			3f��>�.�N��͜>}Z B�;Ｃ�={*66V         ��>����+�eddhĈ.��;<�E������#��Ҍ3���,(�z�.��Ddd�RRRT\\, �����M�F�)         �\o���N�<�peي�n�M���pB�ܹsշo_W
�vxrj��>ӦM����V�Z	���pB˂4p�@w�         �غu�֮]�pe��G��@Ւ�����(�:uJ ��}Ϝ9S��w� �w��N�>�Y�f)\effj��j��7o��a���{Ocǎ         `,_1e��9sF�jذaj۶��ꈈ�Pjj�8  �o͚5.g���- 5G���e˖���@�A�3f�;a�Wj�i�ʕ�ꪫ���!         ��{��U��С����/�&,SA�o���{�1�v@-pj��ɓ�;w��5j�\
�@h��w�yG>��         ގ?�ٳg+\���h���.k��
 ��۷O}��$ 5C���E����D�w���ر��K�d]_|�6o���        �0g健��
G��k����X5���& ���w�u�;~. 5C��&�xY�=����ꫯ�qqq���WYY� ���3g�G��         Li�ҥ
WC�UFF��ڠ4=ǎӂ4j�(�>�@5͛7O���
7��������&d܁Д����?�\ݺu         "UTT(eff���w��Y�w��_W� 	�@���D�S9��֎�t���m����{g���1{k���tvg����*�(g-�H�� B!�����QAr�|>���gƙ�`5\��}]������~7��J=E&���@q����?�|6hx8wxW�^�w�y'�(��>��Ciƌq��� ��W^�e˖��     P2ǎ�ݻwGM�0!~��_e���J(�ڵkǝ;w�w��]��?�c G���C�&S6�gώ���C͕ZPlgϞ���?֬Y      ��o���N����~����RS!p��ٹsg���K1gΜ ������˗c���Q6�Dq�|UWW���� ���W_�U�V�P     P���q���(����X�hQ�PH�{�(�t ����}�˿�K �L�����_����(��>����w(�.Į]�b���     @��h/Mo/�����я~0T��ڻwo=z4�~�� ����ƕ+WJ9�=��)p��2eʔ����;w�P\���Z6ŽR�      ŕ�:u*�&}����,�������Pl���J���k _O�_����6_55^>��,�8��O(�s��ef��     �b���W_}5�h͚51����$p�b;|�ptvv�ҥK�j
V�
iz��mۢl֮]O>�d�pK2�;����x��gMq     (��۷���ts��/�0�cܸqq��� ��w��],Y�DK_C�_�7�(������x�F��Pi��|+W�      �%Mo�ӟ�e��ğ���Y�C-�|555eߵ�t���طo_,[�,���|��g������8Ə0�P�И�     �xv��.\��Y�bE<����%5w(�W_}5���Lq�� p�ظqc���D�̟??/^0R�P'N��ĢE�     �b(�������������&�Ŗ��wvvf�;�ew�O
�7m�eR[[?��OFRڌ�����_�pS�     P;w����G����?������dh �����X�t�)�� w���͛��>�2����S�NI�`Ŕ)S�ʕ+����>�;wn      �oiz�믿e�`��X�xq�p�C9��b���Y�|���{�nlذ!ʤ��1�{ѐ��ܡ<�|������       ����?ǅ�L��4�FB�)�D���� �����@���X�bۗ^z)ۄ�h�1cF9r$�rؽ{wtuu�6      �si�Q�|��ߏ�S�����L�<9�^�@�>|8�=O?�t ��� o��V���ٳcٲe�%�8�#]U��;�į~��       �����O��2I�m�;�	Iip����7ވ���sw��)�'ND�����mv��S��|�}����O~�Ǐ      �'Exe��ߪ��Y1�RSq�ȑ �o�޽q���hii	�+/�6n�e�dɒ�;wn�h�C�tww�����?�a      �/ip�C��L/^���#-� �C�������#p��_��gϞ=Q�����/��I�&E}}}ܺu+��x뭷�^p�     @���O�2I}�K/�0�ry����?�yL�:5 �;dRhw���(��k�:�ɘ�6d�O��<.\�}�Q���      �p�ҥ����L�{�9}�F���ŷ�~;~��_ p����m۶EY�i��?�|�X!p�rz�w�      9�q����닲H7��{�-QWW===���͛�'?�I�g�N�N��ڵ+�_�e��/d�;�NC9uvvFWW��      ����.�����_2������_(��7o���۳��N�N�	�e1mڴX�jU�X"n�r���-[��/~�      `lۺukܺu+ʢ��9�/_0ښ���P2�Ɣ��Q�T�L�N��9s&�=e���?�����;�W
�_~�娩�$     ���2L^z饨��
m�
(�.Dggg�������R{��w�,��������f�ԩY����@�\�~=����v     �1l߾}q���(��s��3�<0ܡ��z�-�;�'p��zzzb�ΝQiz��ŌE��2E�/^�|Ҵ�;     �صiӦ(�4��
�;������I����e%p��v�����Q)6���,m��PN����Ϙ1#      [._��Eve�hѢ�3gN�X1mڴlp`___ ����[�l�_��e%p���m�eaz;c]
[?��� �'mʶo�?���     ��%��[���R��/�0������ɓ�ʕ+��֭[�?�i�������R���#G�DL�2��vƼ��� �+:{���     Cz{{K5<pɒ%1k֬��f���w(�7n�|k֬	(#�;��N7���e���WWW�ei3�W�0�����x��      `lHQݵkע����W�X���ÇP>�������S:)l߱cG�A��h���c]ڌ��r���t�L�     0v���,���b�̙c���P^�p˹s�b���e#p�t8�/_�20����������Ҝ��lϞ=q��͘0aB      0����J31���*~���Uw(�m۶ů~�����S:;w�2H��;::�"m��P^w���"��{.      ]��ݲ���n3�555P^;v�_���R:wJe �+�u��yS#W�ǎ���{�=�;     �(Ka{������n�X6iҤ����[�nP>i`�}�b���e"p�T���[��޸q�bŊy�D<p����z�jL�2%      �;�˗/G̟??ZZZƺ4��̙3�Ӷm���RI�aˠ��#Ə�'w MٵkW���     ��غuk����?����Cy���i�{ccc@Y�)��7ofWu]�R�5k���H��}�;     �(���={�D<��1w�܀<�T@�����)(�;���Dooo]�>ˢ�<jhh�������	���?/^�3f      #k���q�Ν(��}�{y���@����{wJE�Ni�ڵ+�`ݺuy�nH��g�Pn����G     ��J�\L�<9�y晀�0�8q�D�?>fΜPwJ�֭[q���(�����Uڐ	��;     �Ȼ~�z)ڊd͚5QUU�ӦM����{�n �������/�PwJa�޽���E���|'��y��1��<y2.]��=     �������E����Ɗ+�$��S�LɾG�K�N��)�4	����룽�= ��@���{��_|1      )p/�e˖ń	�&5w(�O>�$N�:O>�d@�	�)�۷o������V�\�ƍ�3�;0 N�     �������2X�fM@�������۟��g�;� p����ۗE�E�����S�N�555EUUU)����ѣG�ڵk���      �4|(ݲ[tO=�T̚5+ �RS�k׮��/Ptw
��?�2x��c۶m����W��!#����c�ԩ���P?����w�      �>� ���v�,MpH���>}:�̙Pdw
-�q���Q===�	�����ĳ�>���Q[[�iC&p�;     ��z�j?~<�.��p�����+w�N�N�;v,�_�et����Y�~},]�4֮]���c]ڐ<x0 ���w��qP     `���i�`ѭ^�:�U�j	�s��� �-����Pdw
-M~-����/LuO�{[[�Mc����t3ɡC���Z      �4��*�J,^�8 �RSq�ԩ �����q�ܹ�={v@Q	�)��{��K�_y�l�{GGG<��1u�Ԁ�D���	�     �Ǎ7�ȑ#QtiB���ۿ��V���5 ����t���"�SX�/_����/����-[b�֭1o޼l�N*WUU�6�;0X
�����>      z��틾��(�������̞3f���˳^���> /��� I=ŏ�〢�SX����^:�|�ر�ihh�6o�W��ɓ'�����ĉ��>�����p�B477      Ck�޽QF/^�6��͛���-k%f͚0�8~�x\�v-�H�Na}����û~�z6�}۶m��SOźu�b��Q�TFZڐ	܁�=]�     0��޽[�����'v�ڕ=---�D�����������4�6����s����BJ/�]�zl`���i�b�ʕ�bŊl�6���!;y�d $����     ��9|�pܼy3���ٳٳ~��X�ti6pƌc�ԩS���:;���G	�),�;�t�ԩl"9�����ٕ\�6m��f'��͛g�;�Ήc`���h�5      ��{�_��ݝMt߽{w�H�VbѢE��bL����V^�x1 ������QS#�x�TSH酛���;;;�'������>`8܁�҇��V����      `h�۷/�j���q�ر�ihh��˗��իc����)5w I=ő#G��XP4w
����������T��k�ƓO>0������5�;     �иt�R�?>x8ׯ_�-[��֭[����֭�D�R	iMMM0��?�SHw
'M?z�h0�Ouoii�&�/[�,ƍ�L����q�Ν H</��r      ���p!���ӦM��+Wfτ	F����`�=������F�N�?~\;�Ξ=�=o��f���Ś5kb�̙�V:�N��'�����/      <�4��s���ذaClڴ).\�t#1#A�v���즑����"�S8�FGOOO�ڵ+{�������V҆L�Hq�ɓ'c���     �������s�����ٙ=3f̈�˗g�D}}}�p�������ի�D�N��ǆ����ׯ��K�ƺu벍<,2�~��     <�S�Nō7��w���l���͛���-�g͚0�Ə�&M����t3�����S(}}}q�ر`�����&��޽;�͛��R^�hQTWW|�;p?��      _��^===Y+�������hoo���ڀ����$p�j���E#p�PN�<�Ռ=�*�t� =�iGGG�Z�*�L�� w�~G���w�:$     �ҭ����g�f����c�ҥ�nݺ�1cF��HME� �+W�DWW�ފB�S()|c�K'H�l�[�n��T�ŋGUUU��tڸR�d�# �4��̙31w��      �����i+FIؘ&��޽���ĢE�w�[��Kؼ6P$w
%M'?Ouoll̮�Z�fM�א�f�<yr\�z5 ���;     ��s�ԩ,�f�n%b���z����qxX"V�~���{.�(���=��]��Mu߾}{vB9�TN'��o�+m���`Ǐ����     ��K�];�_���[�n��u��ł�|���� �{<E#p�0>��Ӹr�J�ow�ލ����I��+V�ʕ+c	A����ȑ#0 �      |;i�+c���ӦM�:��KL�81�A�N�555��� IWWW�O��(�;�az{�\�t)6l��6m��fS�[[[��p�p��/f�,�u�      <�Q06�]�|Y+�7JS��a�.��t�m͚5E p�0Lt-�t�t`�{
�;::�\}}}Plw�~�������      <�s���͛7�|�J�M�υ���ѣw
C�Na�8q"(�t���I�K�ƺu�b���A1	܁I��w     �Gcp`~��7o����X�zu̚5+(7Mp?�����BH�\O�>�G:���fOKKKvJyٲe1nܸ�8&M���>�u�V �     ��Do�����v�ʞ�V"����ʧ��) ;s�Lܾ}[CG!�)�K�.�F��Ξ=�=�ׯϦ��kVfΜC:q,f;u�T      �h�;���ĺu�bƌAy�����ݻYS1�����SB7���n'�H����իq�ڵhll      �Y�>�ܹsA���w�y��e�ĢE����:(��ST*������@���"�S�W�7pRyÆ�|��X�vmL�:5�Wj���Z�dI      ��N�<}}}Aq��9E��ihh�Z�U�VŔ)S�b����I�&����`�����@�N!���W�u�V�ر#v���rN�Bx�t�M�     �pR�Ny��y˖-�u�ֿ��/�����X�w�;0؉'�@�N!���7qR9��f�~��     �����ӦM��+WƊ+b�ĉA1��´f`�˗/Ǎ7� ����g�}�~�i��rR9_�N�555��� ��      �� R�aÆشiS,\�0k%Z[[�|kjj
���9s&-Z�gwr��ٳ����ʍ���I�իW;�<Ƥ�)r�x�b �p�B���9�     �zzz��V I��:;;�'M�����b���� �C���:uJ�N�	�ɽs��<�k׮e��7oޜ����[��^�T�ї6dw`���[� v֬Y     �WK��� 8�_WWW6�=�mmm�P@߿��x7�Pwr�w��ݻw�zR9]�bŊl���	��cC<HZ��     ����&i���]�����%
��������6y���ӝ;w`��~�@�N���p�t�RvR9Mv_�pa��kmmF��xk      �o&r�Q�!S�Y�~},]�4֭[3f�ƦJ��p��O`���糃/*�gwrO��p�����T��i[�jU6�}ܸq���b      ��R�����;��{��7o^6pѢEQ]]�-�������e�s��	�+�;�v�֭���OF�ŋ��c���[����W��Y�f�+m�ҩ����  p     �z�;V�+�#�;v,{b����`�)S�c������nw�L�N�]�p!`4���d'����Ғ�Tnoow��0����6�׮]���Q�@-�     �ˮ\����p���زeKlݺ��S�/^UUU��ijj
��H�	�ɵ��hK��ҳaÆ����6pN��t]N�s��<�A�a��!Zccc      �e�6����ӦM��+WƊ+b�ĉ��Ө ��"���	�%������cǎ��SOeWr-Z�(�����w�������ȑ#�f8� _%��      &pg�]�|9�iӦX�pa6���59i�{��:< `@�	��5��҆�����3iҤ�r��M�2%x����СC�k׮8z�hܽ{7 F
��ϟ      |�魌�������̞4Q���#k%����5nܸl(ا�~ ����Ν;Q[[�GwrM��Xw�ƍؼyslٲ%0�T�DUUUY���Ķm۲S� ��Z      ૝?>`���2MuO�D[[[�^�:f͚�t�@���ח5---y$p'�Dm�E�P~����<yr�\�2{�����7n�+W���e-      ���m�0Zzzz����3gΜl(�ҥK��F�6�nݺ�Mq�_Z��+�r+]m��!y�~n�~��x��wc�ٕ\���Q�T�Ҥ��^{-�= ��ҥK     ��������c��ӧ��7ވ���,v�6mZ��]�G��cǎe�N�S�WqЍ<��[W�^ͦbC^ݽ{7��ߟ=iӖ&��X�"&N�E��fq��۷`(�     ���M��
ƚ�7oƶm�b����0����UUU�WK��޽{㣏>�S�N��<������[i
4E�yްaClڴ)�,Y�Mu�;wnE�q��C�ٳ' �R�F�UWW      �3���,�����466fCӓ���ݸq#;�{������G!p'��䖉�Q
�Ӊ��477g'����c���W�������Z,����חE�/     �"Qyq�ڵl �ﾛMsO�D��^�T��zzzb˖-�s��lz;���y&p'�Lp������_�7�|3�����i�'ׯ_����������pIk�;     �	�ɛ4���?Ξ��_��bŊ�8qb�ɡC���^�}<�4D��ݻQ]]�7wr�w�"Mu���̞����r[[[�7.Ʋ������?����:     �e�g��wÆ�d��|Tw�܉�7Ǝ;`(��C���>}z@��ɭ�W���ٳg����}6ս��=�ݛ��c��y�f�����^k      �L�N
8s�̬�H�D]]]ɥK��׿�utuu�P��Wwr�ڵke�����^�����r����֎�?Z����o~�p�B ��tc      _dHEs���x�ײ��˖-�b�Y�fEޝ8q"����;nݺ Ć7�J�Nn	��4�==�ׯ��K��ڵkGu���o�G�	��bM      �E)�M�Ӡ�zzz���s�����������?��?q�Ν w�J�Nn��
_�>�صkW�<��Y�hѢ�����C���͛`$Y      |�����P��7FGGG�755E<x0���޽ �Ś����K)�}�v v�ԩ�ihh�+Vd�ɓ'���駟�+�����0�Lp     �"�Z)��7oƶm۲g��>�3g�������ہa'p'���I��pҟ�w�}7��>o޼,t_�xqTUU����?�1��`�Y      |QPe50���1V�\�=�Ǌ����Wܹs' ��իW�H�N.	��Ѥ��ǎ˞4�}���z��!��~�ȑ8p�@ ���.H�s�J%      p.$����M��w����+Ml��o~c� 0b�	�+�;�t�ƍ ���nٲ%��k��ٵ\i#�m�����lz;�hIuwwG}}}      `p 6x(�iӲ��+V���'��?��������0R$����͛7x<}}}q����ijj�U�Ve��'L��H��֭[�ҥK0���@�     p�i��`�/_�6d��.\�Mu�����СC�s�� Iih`j*F�P<�;��Z)P�7b�ƍ�������۷�h�6      ����^�����3{fΜ�loo����a��������o�)� #-Mq��7wr�w�7pӧO����,v������~tww�h�6      �\
ـ�s���x�ײ��mmm�z��5k֐�o����4�Q����7�;�dJ+�����^˵t��X�n]̞=���{���������A      ��ãK���ڵ+{ZZZ���i�{mm�c��.\�~M��b]@	��%��4���?̞�ܲe�b߾}���k     �����ٳg�g����P��k�Fss���^�������b]@	��%�at����x�k     �{��t#7��������w����X�jU,\�0���������ĉ0���:�\�}�v �'m� �k     �{Dl0������ѣ�3iҤ����b�)S�|�߷u�� m��GwrI� v�Ν      @���ƍ�e˖,^�7o^<�쳱x��/Mu?y�d�9s& F�g�}�7wrI� fm      p��FF��~�ر�6mZ�\�2V�X'N���m۶�X`�;y$p'�Dl �`�      ���`�]�|96l��6m�%K�Ă�СC08�F	�ɥ;w� � k     �{�������w���+��#�;�dJ+ 0��     �=�7 �6 ���R:� 0�w     �{Dl �`����\��� ��      ��� ����#�;�$b �6      ��ͷ �`w�H�N.�� ���      �� �Y�GwrI� fm      p�� ���7����R����\� �Y      �s���  ����UTWW���\J/�  �      ��� �������K��; 0�5Z      ����Y�7wrI� VUU      � �/�{�n@��ɥ�ِ �      ��) ��(L���% 0��     �=w �~&��7wrI� fm      p�	� ���#o�䒈 ��      ��J�  ��*��;�T]]  �      �� ��> o��RM�] �s���     �� �2��F%L.�7.  X      �S�T `0�;y#p'�Dl �`�      �TWW �`����\� �Y      �cB+ p?7��7wrI� V[[      ��
 |Q�ۭ��;�$p �6      ��`  `������;�TWW  �      �1 �ڀ<��K&L ��      ��� &p'��䒈 ��      � 0��y$p'���� `��     � 0��y$p'�� �`w     �{Dl �`���y#p'�&N�  ~     �g��� 0@SA	��%/� �`&�     ��{ `0k�H�N.544 @�����X�     $"6 `0��#%����  �u     ��� �`����\�4iRT*���� ���      �3� L�N	�ɥ���,r�~�z  ����      �SWW�u}}} ��y$p'�R�&p Lp     �\�R�&�޸q#  Lp'���V��Ξ= @���     �E���; �H	��-/� @bM      �E)p?w�\  H	�ɭ�S� ��i�     �� �. ��䖘 H�	      �H� $UUU1a����[&� �5     �544 @:�V�T�F�Nn��
 ���9i     p��ġ7�J�Nn��
 8�     �e�'O  k�J�NnM�81jkk�Ν; ���     �� ]y%p'�*�JL�>=Ν; @9��       _$f ���+�;�6c��; �XZ      �E&L�������	 ��z#���Zsss  �e-      �`ib�'�| @y	��+�;�fj+ ���      ��	� �;y%p'�Dm P^�J�Z      �+� ��RW1eʔ�<��k��� �Sڄ���      _6}��  �+u552a��O.���Ԕ� ��� P.��     |5C�ܬ�3�;�VUU���={6 �riii	      ̰  (7�;y&p'�R�&p��={v      �`3g� ��v#��䞸 ��w     ��6~��hhh��ׯ P>w�L�N�	����      �^
�� PNw�L�N��
 �3iҤl�      _m֬Yq�ر  ʥR�Dsss@^	�ɽ�"\SS��� ��n      �,� @�455E]]]@^	�ɽ���lCv�̙  �aΜ9     �כ={v  �c@�	�)�'�|R� %��O      _ϭ� PN� ���B0� �%n     ��555E]]]��� P&��ww
A� �QSS�f�
      �^�RɾW9y�d  �!p'��B���6e��� [�F+E�      |��	��<RK)p'�AB�Nkƌq�  �-l     ���Vv�� @9477gM%���;w�� J��'�      ��V �\��Ƽy����� ��Z[[     ����J���� ���"�Sb7 (�q���O<      <����GSSStuu P|w�@�Na�嚚���� ���ΝUUU     ��KS�� Pw�@�Na��=mȎ; @1��     �ѥ�b��� ��ɓ���1 ��ʼy�� P`�     �G�n� �逸�
(�;�"z�b�^     ���w,�J%��� (.]E!p�P�y�  ����9�L�      <�����5kV�;w. ��jmm(�;�2y��,~�p�B  Ų`��      ��I]� P\UUU��SO����I�� ��M-      �^
ܷm� @1���D]]]@�)��oݺ5 �b1�     ��kmm ����S$w
�tW (��S�FSSS      ����Ǐ����  �'��E!p�pR�6mڴ�|�r  ��      �㩪����~::;; (mE"p��-Z۶m �/^      <�����N�ӧO(
�;��d��; H:�     ��1� ��{<E#p��Ҕ�J���� �[KKKv�     ��3w��7n\ܾ}; ��H��@��)�I�&�O<�O�  ���,      <����hmm� P&�S4w
+Mq�@���t      �F��*p��hll����"�SXi��o� @~�)"��     :i�Ы�� @1���J�P$w
+�p�Ǐ����  �)�����      Cc޼yQ__�n�
  ��0`(�;��&���I|�A  ��lٲ      `�TUU�cϞ= �[�ܞ:I(�;���8�; ��     `�N� �����'O(�;���ޞ�P���  _fϞ���     ��Z�dI  �gz;E%p��b�ܹq�ĉ  ���v     �ᑆ555ťK� �/��(*�;���8�; ��     `���b6m� @>�7.�y晀"�Sx�ꫯ �'N����      ã��]� 9�x�⨭�("�;���O�̙3���� �C:�VUU      �����㣻�; ��I��@Q	�)�ɽ�� ��ʕ+     ��SSS�-�={� �/�JE�N�	�)��	� &L��}�
     ��Ja�� �gΜ91eʔ���S
s�΍����t�R  c[{{{61     ���4���? ��0���SQ
i3���7n `lK7�      0�&O���͋cǎ �+V�(2�;����
�`�?~|,Y�$      i��� �c���1gΜ�"�S����{WWW  cS� ���6      �����������;���?��a���c AD���QA0"���hS��[�&�$�MbV�ny$�dc��^+I���w<QO0FQ��>_�嚣g���z����-���3���TUU ��Ұ_h��䍂��2dH�q� 䦡C�      ��u�����_= �ܗ6�AC'p'�TTT� G�h�">�O�  n�IDAT��      �v�PN� ����,�t���	��+:t�N�:Ŋ+ �-餕���      �v80n��  r[ڔVPP��	��;C��@J�;      ��}��@=p衇��;y'�i��m� ��ڵ�8       �@nkݺ����!p'�EϞ=c��� ��Ç;B     �����o����  rOEE����!p'/��N� �!]|6,      �;i`��K�.  �2$ _��K�f͚���� �[�{��~`
     @�JS�� �{:u�;v�w�RqqqvQv�=� P���*      Խ�����Ɩ-[ ����o���	��n���f'�      P���n���O>�d  ���� ***����եK��ܹs,_�< ��1lذ(*�      W���w ��{������|�&"�~��q�u� P7F�      �C9$��g�x�� �{i���;y-�q�7Ć �]tPt��1      ����YO�hѢ  �Viii���? ���k%%%1lذ��{ �]GqD      �{�)�w �{C�����|#p'�5J� ��E�1`��       ��������J  ug����H�N��СCx���lٲ  jǈ#���GQ     �\UYY)p�:Թs������בG)p�ZRXX��@     ��5t�����~�ׯ ���5* _	��4(��w�x�w �Y�}�M�6     @�*..�aÆ�]w� @�jڴi2$ _	�!>�$�v;���� �f�3&      �}GqD�}��QUU @�I��JJJ���Oeee�v�m�q��  jF�.]�[�n     @�k߾}���#�,Y @�9������O�f͢��"���  j�رc     ��#Mq�@�I��:v�����	�G������Z P���bРA     @��~��~ϳf͚  j^�!�	��:t��rH<��� T���:*5j      ����1jԨ��� �Y�[���;�;��c�9F� լY�f1r��      ��9������o��7 Ps�<��ls�;�;��8 z��K�. �z��&M�      �OfTQQ��{o  5���$F���vh���w �&���ٱ�      �_GuT�w�}QUU @�>|x�������7:w�˗/ `�92Z�l      �_���ѻw�x�� �^1z�� >"p�Hocǎ�+��2 �=רQ�l�      �߸q�� P�ڵ�#w�C���n�-�z�  �̰aâM�6     @�׳g��֭[���� T�����ww����q�1��UW] ��K�G}t      �p�;6.��  �G�^��K�.�����СC���o7� �@����,     ��e���ѡC�x��7 �{���g	���ɳ&L����: �]gz;     @�TPP�Mq��/~ ���ܹs���3�O��NTTT�w�a�; �4����<      hxRKq�-�Ě5k �s�sL�y�4�;�D�@��D���  v�Q�F�{'      SQQQv����  �Lǎc���|��vA�y��?�!V�X �9rd�m�6      h��������w �C�&M2�>��vAz�<yr\r�% |����0aB      а�)��Ǐ����7 �:��_@�����ѽ{�x饗 رѣGGYYY      ��UVVƝw�i�; �c�=��v�w�S�N���� |VӦM�)      �S�`�u��1����n�ѣG���;/^ ���7.JKK     ��������U�V �s�'O6�vB����㏏^x!�m� �GZ�jGuT      �_���'�5�\ ��ҥK0 �/&p��ԩS�8��� �#S�N�ƍ      �gذa�hѢx��7 �|��0�vN�{�㎋�<6l� ��:w�     @~*,,�ɓ'�e�] �����#z����	�a�l�2Ǝ��rK @��>}���      yn���q��+�� �gM�6-�]#p�=4~������c͚5 �*���gϞ     @~K��L�?�� ���Wt��-�]#p�=T\\�w\\u�U ������b      >֫W��۷o<�� |�Q�F1u�� v���BEEE6�}�ҥ �f�رѮ]�      ��N8�X�xql۶- ��Q�FEyyy �N�{!�5s�̸袋\��W���b	      �Ծ}�9rd�{� ��Y�f1q�� v���R�Ν]��w�O�%%%      �h����裏Ƈ~ ��R�^ZZ���C58���'��>�  ��;��c���      ;ҢE�?~|�t�M ��m۶1jԨ v���A�a5eʔ��� �F���'�      �g�ر����ʕ+ ��	'�EE2]��s��TVV�C=/��R @Cu�QG�~��      �ER�7}����K �M�^������;T�4�v֬Y�����u�� ���u��1q��      �]�¾�}�Ƴ�> �/�&��N:)�='p�j�&ڎ3&-Z �Мx�QRR      ��fΜ/��Blٲ%  �����<�='p�j6iҤx�'bժU š����      ��ڵ�B�;�3 ��kٲes�1��;T�ƍgǋ\|�� AӦMcƌ      {b�ĉ��#�Ě5k ��W4i�$��#p�зoߨ����~8 ���>}z��>      {���$fϞmX  Z�>}bȐ!�=�;Ԑ�3g���?k׮ ��z��#F�      �iX`���㩧�
 hh���㤓N
�zܡ����f��/�� ��h�$����      ���¿_|16l� АL�81ڶm@��CJ;��?�x @}3u�T_      T�����4iR\�� EǎcܸqT�;԰�O>9�,Y��~ @}ѭ[�5jT      @u=zt<��#��k� �w1{��hԨQ �G�5�y��Y�~�e� �%%%1w���"      �Saaa�r�)���~7�l� P���[ݻw�z	ܡ4(F�<�@ @�;��]�v      5�S�Nq��Gǭ�� P_�n�:�L�@��C-�9sf,[�,�z� �\էO�9rd      @M�8qb<������ �71gΜ())	��	ܡ��7�y�������غuk @�i޼y�z��E      Ԥ���8�S������z���2z��@��C-�ҥK{�q��7 �Y�fE˖-      jC�Νcܸqq�w �eee1mڴ j��j��G�/��K� �#FĠA�      jӤI���矏W_}5  ���ٳ�iӦ��;Բt�ּy��_��_b��� u�]�v1cƌ      ��֨Q�8��S㢋.�M�6 �ѣGG߾}�Yw�鈒�����/ �KEEE1��hҤI      @]�СC����_�:  W����S�P��PG��� ԕ�ӧG�Ν      �ҨQ�b�����SO �����đ��� j����I'�˖-�իW ԶtdV�A!      �9s�ī����^ @.�4iRt��5��!p�:Դi�8����G?�Qlٲ% ����q�i�EAAA      @.hѢE6��?�iTUU �=z��G@��C�֭[�p�	��_�: �64j�(�`UZZ      �Kz��Gyd�u�] u�Y�f1w��(,,���!�5*^{�x�� jZ�Xս{�      �\t���ǒ%KbŊ u�K_�R�n�:��%p�q��'�o���� PS=��l�      䪢���7o^\t�E�y�� ����0 ��'p�Q\\g�yfvq�� T����3gN      @��رcL�:5~��� Զ�>4}�� ��rH:���N��/�8��� �K�&Mb���-      ��G��%K�ēO> P[JJJb�����Z�n�!����'&O�7�|s @u(((�SN9%�]      �E�=�ܹs�{��^��� ���O�:Pw&L����z��/	 �['N���      �7���:+.��ذaC @M:��#cذa�-�;䠴��SO����ov �W����{l      @}U^^�Mr���UUU 5�k׮1}�� ��rTځ�`����w�k2 {$����N�6N     @}6`��;vl,Z�( ��5k�,�8�(*��B.�9�}���$��.��d vKiii�}��Ѵi�      ��`�ԩ�bŊX�xq @uI��͛mڴ	 7�!�80�L�7�tS ��hԨQ̟??��      Eaaa�~�������z�� ��0mڴ�۷o �C����	����/ `gN<���ٳg      @C�N2NÞ~��Ė-[ ��СCcܸq��;�'�tR�\�2^|�� ��3~��8���      ��]�fC����� �=թS��3gN �G��D�F���3ό�}�{Y� �h���1u��      �����2^y�x�� vW�-b�Ѹq� r���t��W������k׮ �.M��;wn      �Y�f��o�K�,	 �Ui��g��[� 7	ܡ�iӦM�s�9��(6n� жm�콡��$       _�@q����}/V�\ �3ip�)��|p �K��P�.]�d�\rIl۶- �_�Ȭ/���-      ����8������~�_�> ��L�0!�@n�C=u�!�dGm�� �S�ƍc�Ѯ]�      �|վ}�8묳�'?�Ilٲ% `G�'O �	ܡ9rd�Y�&n���  �řg�ݺu      �wtP̜93��� �t��i���>�;�s�&M�M�6ŢE���PXX��zj���7      ��~����;��w� �]۶mc�Q\\@� p�`ڴi�aÆ���{��-�$�5kV2$      �O�2eJ���{��� 4o�<�=��hٲe ����;�|�ɱq��x����k���1r��       >+5�g��"��{. �_ib��g�����/wh �ک��[�n��{, hx�N�GuT       ��Q�F1����˗/ �Oaaa�~��ѭ[� ��;4 �My�ܹ�$�g�y& h8�=��8��      ع&M�Ĺ瞛E�+W� ����<@�$p����(�<����OK�,	 �ѣGǤI�      �u��O|��_����z��  ?��1bĈ �/�;4@���q�9�d���e���k���1cƌ       v_YYY�w�y�$���{/ h؎;�;vl �������,r�����믿 �?��9s�dGg      {�]�vG��֭ ���:*&L�@�'p��iӦ��/9~��śo� �)n?�3���0      ��ӱc�8���A��ׯ �#�<2N8� �;4p-Z��o|���$^}��  �2$N;�4q;      T�Ν;ǹ�?��c�ƍ@�p�a��̙3h8��5k��u���K/� ���ʘ5kV      P��u�.����g�y�� �~4hP�r�):h`��}۶mU4hM�6��|�+q饗���? �Q�Fŉ'��      jPϞ=�3Έ�.�,�n� �O}��y��Eaaa ���}[ ^III�s�9q�WēO> ����Ǵi�      �y�����O?=k(�S �Oڬt�YgEQQQ O��]����=�B���+��� �V�֞��q��      P{_�җ�k���#|p,\�0���h���>�AI�{څ�&�?���@�Hq��3b���      ԾaÆEӦM���/�-[� ��o߾�`�q;4pY�m�6�!��)���]���O
 jWz�3gN><      ��ӿ�8묳��?�yl޼9 �M��z���ـW�a����yh���&M��m�� Ԏt�5o޼��C      ��_�������cÆ@n:th̝;7(4|Y�y�f��@�<yr���č7�UUt �IiSQ�MܧO�       r�A�~���?�u�� ������O>9�
�,pߴi�������m۶q�W:n���l�2�9��ҥK       ��k׮Y�����$��� �n��m�ԩ�v�3Y�q�F5+��V�Z�%�\�"���k�.�=���      �]�;w�����o��o��� u#��ӦM �l��.p2ݺu�/�0.������� ��ںp��hѢE       ��}��q�d���U��ړ����1v�� �S�oذaK ��6m��7��l���e��=7x���;wn      P�~�k_�Z��\�2 �y)n�5kVTVV����}�ƍ&��RZZ�~�����~8 �}�G��3fd_      @����ƅ^�^zi,]�4 �9EEE��C=4�������� ��?0�m�6n��� `פ��ٳg�a�      @����w�yq��Wǣ�> T�f͚��G��=p� ;��O�4)Z�n�^{mlݺ5 �|�[,��:(      ��!��7o^���P�R�v��F� ��w�}wc |��ÇGYYY\q��nݺ �:v��&N'_       ��!����կ~eH @5�o����=��l�}����Q�F�yz����ַ��K/�7�x# ��~���i��M�6      ��9rd�j�*.���ظ�\Q�=շo�8�3�I�&�IE��|��Ѽy� �"i*�7��͸���'��|��4�7.�N���      �e�~��/�5k� ����2N>��(,,��q�~�z�;�KJJJb����hѢ������* �Q�A<w��0`@       �e����/�0~���������KA��3��#����q�nݺ �UiJ���㳋�+���k�w:v�,����       �S�V��.�+��"�y� ��A���~zr�!�E>�׮] �+����|'.���x�� TTTĬY��-      ���~o�p�¸���㮻�
 >+<묳�C��3w`�����׾����\�ZQQQL�6-ƌ       ��̙3��_���y�� �#i��y�Y�f�+>���� �S)��~�v���ƍ�!�w�}c�����      ��:4�N|饗��ի �ĸq�b�ԩ�}�]e�;P�҅Z�.]�+���˗@C0p��8�S�$      v�s���o}+.���X�dI 䣒��8��ScРA���@�+//�/�0n�ᆸ���* ����l�1c      `W�h�"�?���馛bѢE�	 ��~��3ό���/ ��ǁ�{� ե��(fΜ�rH\u�U6� �N:6��3�p�      ���6mZt��-���X�~} 4t�/}�KѴi� �S�k֬	��ֻw��������+��_�\WPP�F���?>��      �7�غ���cŊ��M=�w\�?> �ƺu�����m۶�E�:�j�*;v���������iӦ �E-[��9s�D�~�      ������7��͸��⡇
���u��1���ڵk �w�y���֭[c�ڵY�
P��D����8���i�z �A�ŬY��y��      P�7ns���n�򗿌?�0 껁f�KKK�:|*p�����I�ȭ/�0n���l��# �R�&Mb����&      ��6x��l������/� �QqqqL�:5ƌ �i͚5��� 5�Q�F1iҤ�ݻw\s�5��[o@]H�Ci���       ��u��q��m�ݖ���� �/Ґ��O?=:u� ��3�W�^ ��{����|'n�����`�;Pk�6m�|�92


      ��f8��l@�ڵk ����#���ӧg�j�g�U�V@mJt�M�C��.֖/_ 5�o߾1{��(++      ���~������q�u��_�� �E-[��9s�D�~��&���۟�W�\ u�s��q�f�n�y睱u�� �N͛7��3g�СC       ��h�",X�?�x\{�~�� ��ʆ	���@MK=���EEE1eʔ6lX��W��^x! �V:���";+�P       W<8�v�W_}u,Y�$ �R�&M�ޢ��2 júu벍~�
��y�زeK�ԕ���8�����믿>>��� ��ڵ��O>9z��       �A�֭�_�j�u�]q�M7ŦM������7��^VV �����n?U�WUUŪU��}��P����4ɽw��q�7d�{z���5���:*&O�l�      P�nb̘1ѿ���//��B Ԇf͚Ŵi�Lm��ʕ+�ۢ}A�䊖-[�ܹscĈ���&�x� �"iZ�̙3�C�      P��i�&�;Ｘ����w��]lذ! jJ�~�b֬YѪU� ������ً@.9蠃����v�}��q�-�ć~ �Զmۘ:uj<8       �4�=MR�ӧO\w�u���@uJCH�0�C=4 �R�ؓ����_ f�o6,n���,v���
 �5n�8ƍG}t      @C���ƹ�O?�t��W��5k���Hh***bƌQZZ um{Ǿ�	� �,}�J;��_}������Y�w\���      @>�ׯ_���#���+��ضm[ ����/f͚ݻw�\�>Ӭ\�2����=MDN�@.�֭[|���v&�������~;������O��"      �KM�6�x8�u�]+V��]Ѹq�8qb�;65j �⭷ފ-[�d�?�oڴ)V�^mڴ	�� �L�ӧO�+��[o�����0�k�.��>h� ��      �����}��ߎ�~8������������O�֭[@�ICڷ+����׿
܁z%�&3fLTTT�����{ol޼9���e˖q�1�Deee       I����rH60ܶm[ lW^^�������ԯo��B���_�v� �7͛7�3fdG��v�m���h�z���$F����M�4	       v���4X;���o~/��R �-u���0a���@�[�|����v������,fϞ�}@K��Q\UUU��*��eʔ)ѢE�       `����q��O<����cժU�t�CEEE��Ѳe� �Ҁ���@���י;wn�3&;��駟�C+..����?~|�j�*       �})n<xp���/��l8��h�z��ӧO�N�:@}�~��X�f���a�z������y������.�7�x#n��l���r�����{��      ���!ci�؈#�^�{�m۶��t��!��~�!�@}�����,��'�)�i'@C��~������}ѢE���ݡ	�      j^t:s��8�����o�'�|R/D�֭cҤIQQQ���P����>7pOO�U
��Ν��R���;��G��[�P;�4iÇϾ��       �#Mx^�`A����D���~:��)m\7n\�=:;��>K��?�s�W^y% ��;f���ɓ��c<���q�� jF˖-�� cƌ�f͚       ��k׮q��gǲe�⦛n��K�P?���ĨQ��c��4/����,p����IGqM�81����{�>�z�o�>ƎÆ����       ��x�����=���,tO�݁ܔb�#�8"�>�hC����ߏU�V}��-��}��X�fM���@�HG�L�4)&L��=�X,Z�(�x� �L��ݳi�����        ����+[)t���G�"l��ޞ|��� �&M�N���J�q�u�]��%�m��K�?�zh�7.��o�       �~��?��q�m��08jGiii�=:,شi� h�v������@�K�q���[o�����ğ���X�~} �ֶmۨ���#Fd�!       P?���7[i(��w��<�LTUUP�Z�l�~xu�Q�v /��w >R^^3f̈iӦ�SO=��w_v4䳂���ٳg�80
      ��a�P�+V����x�Gb۶mT�4X��#������� ��s�k����ǿ0pOaӦMѸq� �#EEE��i-_�<���裏Ɔ�ž��Mj9rd�j�*       h�:u�s�΍I�&e������ظqc {�G�ٴ����g���믿�����-[�dS��dV >�s��1{��9sf<����T�^x��\4HisG��6lXv�i�       ��M�6q�I'�ԩS��?��O�z�� v��#��ݺu�|�dɒ>���{�t�R�;�N�c��Ou_�jU�S9-q4]�v��Çǐ!C�Y�f      @~kҤI�3&F��<�L�u�]�����Ś6m�vX�7.��� ߥN}Gv�^������H��^{�x衇����k���[��C=4F����       ���� ��뗭7�|3���l��ƍ��.]�DeeeTTTD�ƍ�����x饗v����Jl޼9�N��IN�:���_�b�'�|26l��kZ�j��N"�޽{��       �:t��3gƔ)S��G�{�'V�X���IC��#�8":w� |�o��֭���v���=E�tP �g
�W�^�J���X��<�z�����J:�o߾�n�t���      ��JQo�T�ֲe�����'�x�Tw�F�n�b���1t��())	 v,�<;ܓb
��G:c��\۶m��_~9��{�X�vm@Mkݺu���ߤv       jԁ��Y�f��O?��w_���QUUА���ƠA�bԨQѩS� `�}�����.�/Ύ��z�i��/�N8�X�|yvA��3��k��Pҿ�t��!��m����E�       Ԛ40aK뭷ފ?�������;�P_e-�a��ݦ>�]�y��X�t��~}���_=֭[��2�f��]�t�֤I�����B���#��:���ݻw���o߾��      �	���q�q�e+�{衇��G���? ץ��ݺu�6kTTTD�������/~a�K���m۲�aҋ2 ��m۶1z��l���?�����q�x�.>i����={F�^�⠃�F�       �� �O��/�Gy$�aÆ�\����]�Ɛ!C��C�}��' �;�>��~}��$E�w�����J�rZ�ڵk?��S��r�� �l�{��E�)h/))	       �o� �tByZi`j"R���O��N�HQ������L��۵k T��{���ˁ{*�Ӵ���@�jٲe��9�$�K�.�b��^zɄ�h{�޽{�8����͚5       hH��~��e��O�_|1�x�,xO}Ԕ��"8p`�Lj�i��Ά��r�f͚X�bE��[R�N��~�F:��W^ɂ����}ݺuA��.��1li7p
�S�޸q�       �|QTT}���V�׿�5�y�xꩧ��_6���VZZ={��xS�a� 5/]ߙ]ܓ��@����4i�M�N+It��߲�=�˗/�6-����6(��״R�~�DYYY        ױc�l�?>�}�ݬgK�\�����LAAA6l�w��YО�� �����sv+pOǼs�1@��>�w��![Ç�K���o����)zO���Z�z��5$�,o׮]v�ݩS���vGZ      ��iժUTVVfk۶mY���/���?K�.�-[�$i�`�=�A�)j�i ԝ͛7ǒ%Kv���
�_}��X�vm��@����[�5x���ߴiS����J�{���B��қ;���j۶m��v�Ƃ��?       P}���Ӊ�i����D�ϥ��˖-������6?t�AY�~��Gyyy ���sjwf��4�7�}�/ O�ƍ?��������J��ʕ+���;�|��{ｼ�,..�����w�}��6m�|����͛       P7�4i�M�N+I��K/��MvOa]
��k8R�ѽ{�����n ���{�]z�n��O<!p�Ci�{���J�(��)rO���5k�����V:�#���׭[~�a��ߗ&��h��㕎�J�z:�$�O;|SԞ�       �)x�ӧO���8��S��&����kٟ��?r[IIIt��)�x��f����xꩧv�y��/^�8�KKK �K�}m�w&]��}����Ziwt:~d�ƍ�u���9�o?i��?)MUOk��7m�4������4�>�O�����o_�b       h�R�бc�lUVVf�}��Y�|��W:�^�^wRϱ���G�Ν���o�>kB ����U�v鹻�����'��#F ���޽YU����c} �����$jlJM|%F�ֶ��M��δ��&M�S'�tҙ���bZQ�5���@�"��G��օ]XvY��.��۞�BMb"�}�{��3�s��=砻�}��ږ�       �PK>���[��\.�x�hjj����ؾ}{zL>Ş��,,L�����~�A��z�@�X�r����������         �����'N��Λ%�ޓ�}ǎ���;w�L��'[i�O�筍;6N?��ÓD�g�}v�v�i�V} J[]]�������ק�B;餓         �E����.H��
�Bttt��{[[[�޽��$�'�8p JQ��|�����$dOfܸq�ׇ���Ç �)�4��MaG��|>�V�W]uU         @����8w�&]]]��ٙ.�ݳgOz<�8�������><�\.�BUUU�=���5*��IB�d���'3lذ ���r�ʣz�1��˗�        �UWW�3~��#z}��P���חｽ��$��e��^��%�9�~��d���M�#G�L��$^O��#F��O��m���t�G������]c��rJ          �+�
h�: ����hii9�s�9pO��UWW�\sM           ��-[���9��=����          �f�B�+V�y��oڴ)v���ƍ           H�_�>:::����
ܓ�>��~���           $�.]zL�W��X�xq|������           ���߿?V�\yL�w����7n�.�            (o���ӹ��'�-�w           �,Yr���K�����ԧ>���          @yjll�m۶��������k�?���           �i����u~��E�	�          �TOOO����u�~ܷo�1a           ��$q{.�;�k�[��H���          �Oғ�~ܓ���o�ѣG           ��7ވ����N��i�~��W           �?��'�5pO���+q�UWEEEE           P�zzz����_���{SSS�[�.���           �m�������/����=1o�<�;          @����`��~�ހ�?���c۶mq��           �iŊ�k׮~�ހ�_|1n���           �4͟?�_�7`�����S�L��c�           ����>^��~���}}}��K/�'?��           ��̛7�߯9`�{b��O|"F�           �����X�zu�_w@�\.K�,�뮻.           (s�΍B������=��/Ƶ�^Æ           ��޽{���v@�=��{{{{�X�">��           �m�����; ���=��/�����FEEE           P����.��J���Ԕnq����          ����/FWW׀]P��̙3��.����           ��twwǂ������Ĳe�b���          @q�;wn��A����/�<����           �}���K/�4���Ҽ��-�.]��G          ����s�E.����*�9s���ɓmq          ({��W^yeP�5���ݻc���q�5�           ٖlo?p����kH֨?��q�W�	'�           dS��|ѢE�v�!	������          �lJ��<xp��7$�{��矏�|�#1r��            [v��?��O��C��ݻ7�ܧL�           dˏ~������{Y���7o^\q�q�g           ٰaÆ�����i�~��������o�=           z�|>�z�!����_�n]L�4)           Z�-����!����������          ����3g��3�777��ŋ㪫�
           ���ٳc߾}Cv�L�g�y&>��Fuuu           0�v��/����2�wuuų�>7�|s           0����+�����ߐ��=�`�����?g�uV           08֬Y��P�T�����G?�Q����m           0�����,�T��H��������K          ��5w��رcGdA����?^xa�=:           ���1gΜȊL�QSS����          ��W(������ȊL�ŋ��_]tQ           п�f{����%��������c���          @���쌚��Ț����֘={v�t�M          @�x��ǣ��;�&Ӂ{b�ܹq�e����           �U�VE]]]dQ��|>������O�Æ           �M.���{,�*�{���)�ϟ�_}           pl�~����般*��=1k֬��K�3�           �N}}},^�8��h��������aÆ           G���'}��(
�eE�'�瞋o�1           82�=�X���F�U���3gNL�4)&N�           �v+V�����(E��������_��c�ȑ          �[koo�3fD�(��=�k׮x�'��[o           ~]�PH��wwwG�(��=�t��x�{��Ї          �_6gΜ����bR��{�����'Ʃ��           �-[��g��bSԁ����ӕ�������          P�zzzb������Ŧ��ĦM���矏?��?          �r��ODKKK����gώ/�0&N�           ���W_������bU�{�:ڴiq�=�Ę1c          ���ر#f̘Ŭ$�Dggg<����/|!��J�?          �m�r�tixr,f%U�o޼9jjj�[n	          �rP(�?�Al߾=�]I�����y��'O          �R��s�E]]]����3f̈��>;�=��           (U�֭�Y�fE�(�����7���o�=�����          Pj����{��^���(%�'��~����������          �R�,��w����RR��{bժU1gΜ���          �T<���e˖(5%�'fϞ�x�;��/          �b�p��X�dI�����B|��ߍ��+�=��           (V6l���z*JU��\.=�P��?�c�;6           �MsssL�6-<��,�DGGG<���q��wǨQ�          �X�ٳ'�N����Q��&pO$�X��w�w�ygTVV          @�����q��ݻ�ԕU��X�vm̘1#����<           �,������c۶mQ�.pO,Y�$�<�̸�           ��|�����~�,�ď��3fL����^           d�/�/��r�����B<��q�i��ĉ           +V�\�.�.7e�'z{{�[��V�}��q�g          �Pۼys|���O�z���������/��t�;          �Pijj��z(]�]��>pO������ߟF�cƌ	          �����<�@twwG�����;wƽ�ޛF�'�|r           �C=sggg�3���z��������          �������tttD��������:uj|�󟏑#G          �@ٻwo��{׮]���-���������>��1bD           �����4n߾}{���`���1mڴ��;����&          ���r�4n߶m[���ۿ�������������          p�8���7���1�e��QWWӧO������aÆ          �����I�������	܏�����_�������Ç          ����S�FCCC���Gh�������w�#G�          �#�w��x��b۶m�o&p?
�� �w�}�w�wQ]]           o���3퐛����N�~������}�sq�'          �o��֖�ǭ�������[��׿�����?cƌ	          �_��Ғnnooo����m߾=����������i��           �$�q�����#8r��k׮��7��F�g�qF           lٲ%x�����
����8�޽;��~�w���          @�Z�vm<��Ñ�傣'p�����&��n�->��          P~�,Y�=�X����F��Ozzzbڴiq�-�ĵ�^          @y(
1gΜ�5kVp|��(�����عsg�|��QQQ          @�:x�`���G,[�,8~�0��hkk��n�-N8�           JOWWW|��ߎ�7�C�>@^{���7�w�qG�|��          ��]�v�ԩScǎA��������W�w�yg�?>          �������ַb�޽A����_��W�����.          �x�X�"y�������}tww�}��S�L�n�!          ��R(b�ܹ���8}����|>555�������cĈ          d_WWWL�>=֮],�� [�lY477�����~z           ٵm۶�6mZ�ڵ+x�!�lq�������[�K.	           {jkkcƌq���`p܇H.�K��q����M7�          �|>�<�L�������B���ҿ��q�m���ѣ          :��|'��'pπ5k�Ŀ������g�}v           �o�ƍ���Gggg04����_��W��o�+��2          �������矏Y�f��:����3f�ڵk�3��LTWW          0pv���<�H���CO��Auuu�y����g?_|q           �o�ʕ�ꮮ� ����=�P|���O~�QU�G          �!����O?�-
�E5�a�B!�ϟ�֭��n�-�9�           �]cccL�>=Z[[��������򗿜nr���k���"          �#���c޼y��$����l�����x��'c͚5���~6N9�           �^[[[<��#�q�� ��Ef�ڵ����q�M7ŕW^          �[+
�x��x��#���'p/B]]]1cƌx�������bܸq          �����x��G���>(�"�f͚����������xTVV          �����x��c�̙q�����܋܁���&~����g>�?~|          @9jhhH��777�I�^"6o�_�җ�뮋?��?��*?Z          �C�4z���1o޼���A�RA����^x�X�zu��}	          �l͚5���G[[[P��%(�H��~��q��W��ܫ��          JI{{{<��ӱ|��t�KT�P��_~9�-[���Ǣ�ʏ         �����,�9s�DOOOPZ�%���;jjjbɒ%q�-���_          P�V�Z?�����-(M�2���S�N�I�&ŧ>��?~|          @1غuk<��S�q�Ơ�	��̺u��K_�R\s�5����1jԨ          �,ڷo_<����K/E>�J����������c�ҥq�7��{eee          @$���'?�I�r��|��XWWW<���ӟ�4�L�_|q          �P)
�lٲ�5kV�ܹ3(?wb۶m1u�Ԙ0aB|�������          �%	�W�^�nlojj
ʗ������fL�81��O�4.���          ���nݺ�����[���5�7o�{�7���wŔ)S���~w          @J��g�y&��mڴ)����ǤI�⦛n���??          �x$˘�����>�W	�y[ɻc֯_�^zi���Q�s�9          Gc�ƍ1k֬ذaC�o"p�
�X�re:�z׻�n����}QQQ          �V�u�����s�ECCC���s�6mڔN����k��ɓ'����          ===�lٲ�7o^���)�;Ǭ��)f̘3gΌ���:>�я��ѣ         ��w��X�pa,X� ������������f�J�a��8���7n\          PZ[[��_�W^y%z{{����~���b������/�<����x�;�          ��B��ׯO��5k֤_�����������6��������率�O<��          ���ٳ'�.]�nkߵkW@�3��o�5551s����>W^ye\t�EQQQ          �C��-Z���Z����Aq���X�bE:g�yf����+���N:)          Ȧ��������F[[[�@�3�ZZZlu         Ȩ|>6lH����ե_�`�3d޼�}�رq�e��?���0a��         `
�hhhH��W_}5:;;����Lhoo����3nܸ���K��}�ĉ         @���Ew2g��݇c�SO=5.���;         @?ٲeK��֦a{GGG@��ɴ���ñ�Yg����Ɍ?>          x{ɦ����X�|y����d������ܜάY�����y�{bҤI����7F�          �BWWW�_�>֭[�W�����!p�(%��-Z�NeeeL�0!�����E]�w^TTT         @�H��oݺ�pԾaÆ����F�N�K��nڴ)���'��nwO���8jԨ          (5���KC�$h_�jU�ٳ'��	�)9����t��t�����|g\p���w�;��>bĈ          (6]]]�q�ƨ��O�۶mK7�C)�S�<��O&1lذx�;ޑ��'NL���N:)          ����-bӦMiԾ}�vA;%O�NY���͛7�s�駟�nvOb�d�9�t�;         �`��r�u��4hO���_���΀r����ܹ3��������������8�����Ϗ��ǧ����         �xuww��طlْN���� p�_��磹�9��K�~~̘1i�~�Yg>&��G�          �*	ٓ%�I��t����v�
�	��utt��nݺ��UTT���g���駟�N����N��#G         P�:;;�`=	ٓimm=|ܷo_ GG��!�(����t6l��k�5jT�;6N=���8nܸ�x�'�)��'�tR:Æ          ;8�����ݻ7=&�r������w���� �ϡ�����_VQ���QOOO�ر#�ߦ��:�ޓc��}��ч'��G��F���UUUq�	'�����Ǉ$߷1        �r�,������璖/���������/r�\�'����$�O���+ړ��4;��笇.���{�ox�{��}����* (&�w�u��        8F_��ϫ���@Q�,�l�뮻FE�*            �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��       �v�X    `���4vG   � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �  Ԯ�6 �h ���T���,Sĕu�@�'pg���8        �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��~�y�_˲� �<ϗ       ��^��x <�i�~O��~Ǿ��[>         /c۶�[> ���           $��k����    IEND�B`�PK
     ���Z��n  n  /   images/a46afb92-29a7-4c70-92b4-1e1235f7410a.png�PNG

   IHDR   d   �   +n/�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��io[U��Wl'q�fh�6miZ(P(C�2�|x��
�*\^!U�B|������ $�2�I@�g(3�<�i�$�<��ݿm/�4��Nb;��U�:�9�׸�^۷v�Z	����as�J|*0���o��Y�FNt
��[�1m_��?(}Q>P y�2�I�2��d��0��a�$�(H�Q��< Fy@2��d��0��a�$����SOɓO>)Ӧ�1���/((���By�g�D���!x������<�hKKK�u����TWWK �/�A�_��|�/F#�x�
JKK�D�U�V�=z���s���/���<���E�Ge}��O���.�����r�9�șg�)ӧO�_�F��2�O�W��ϟ�ɕ��Ef@���� '������o�m۶�P�%<���򴵵Y ���3g��2(�P]��G���zc�� ����<>묳���[��w�{�C���t�M�b�
��@;O�!� GU=����7�xþf��E]$w�u��D�y��C��}��7KGG�lذA|xW��8��8r�<��#5��z����_����eƌqՔ�� :88h?��,..��<����ò<`䫗
�U܈�***�ꫯ����� ���#�������r��!�wsB<1<�e˖Y`���O(�Q#�{�n��?d������ky?/^,K�,��<s#@����R,@ ��_��_]�9b_}e:�mٲE>��+v�^{�}�D�xs��ak�qaǒqi�o������n��.���%ڀ�u�A��5��������k�9��ڱc������}�Q�n�:9x�\��8�r����s�=g�ǢE��s���)���q�mmm%��}��ɽ�������NXTT$?������L��>Y�`���w#F�����+	ut��y��g���ώ�/�Ђ�:��h6���>��o=Z7�D����nG<����=�!?L�%}��6�d��ZL�qګ��j���[��K/����!��������vl�駟�7Q�~����|�r����~���	I���g>��SH���x��N;�4��#�@%�p�裏�w��~�Ao
�{@
���ᤵ��V7�L����%����#�i�&�=JJJ����'*͍0�dxq�4���@PI���f����I֯_oG<��t�RkS���c^4�sҪ���u�jµ�`��/�l@E�}��V:b����Μ93> �'F���h�y<b�J�g#�l��Ih
��~+555�����7�6�-k	����u��D�H4¦&��� �JB��ro�n3�%�C��`?�s�o"��ƛ��pR� ����ܹs�n�AG{�z�68�(()�� �� ��_|1a��#%�\�*� �u�1�\`A��W�w�6���'�������/�8���� F�HU�@�͛'W]u���/�]����\S'|�y�g�ډj���ґ�(#��P1�P)�}T���'Su�o�ݺ��[���<`y4��	�0��裏�+��"�y_7"2_�j�̚5+)ҡ �t�v��dp8t^�kU�G�hpL��<���L��c�=&/���͆�#�{T�Xj<f�#�?��CV��k�ڵ블	7���f`w��ɂSQ90~�޽6�RCc#��jj�#Xm���=��q4��xnj#⻤����P�H�XUI��95̡ǳ�q+u4�{�6e���q��o�H�����Ǎm޼�zy���n���M��&���ß�)�g϶G�~s���d2��kll��L��ʄ/'�tR��Od�&\J�?� 8/�c2�����n�߄Yc��t:�q�Pka�atõ��7��T�s�ZhH���x�sq�\+��)��r�{\�x4Ƹk{�m a8*f�ƍ�@j�NrdN�<���eV���5Sf�AQkF^yY��N�F���_::�䰑��C����Ez��#��B�0#Q�ؙ�J�+L�2���E#����Q�,np��`�a���e�YK�43�j���Q������2��2��a^
T�6��J�4̑�b����a���l���wȠyn%J�͇�3~��6͚�L�I�(3��O?ّ�TM#L#�/�@�_|�̬��ζViڹU6:(�248��Q���{
�WX$e�RS7S�<�t�	�ɮ��rd`� � �R���[���Λ�)��7Jf�:$5�j��������/)/.��[7��쐞��F�cm�S��Q� ��~T:����l_(�J�>���A9�;$�<��ະae
 *ݩ���`|��W֋rf����"�,�V"��e���d���� �����{b�|pN{d�%2��H�t�38q a���V���⊈�.J �����TQH��r�,�.�B�G�6J��	�`T'���3�,/�ș�e��{P{�1��T3�H��S}�F�/��b� c4�߂�2i�*������_Zp4@C�_J|���/((OXRv��i#~���	"�Ci��۳g�5�c��)5e2Ϩ��y5*-�J��k������V�l$L�QA�r@{�׿��kk #	?É��K�'a�f��k)���Ԑ�*	��Rm�S7�\<�AUU��܊i�V�`(q]uFR��h��5�H
e�����ȓ�kQ0 �ʸ���L,5���I�p@Z��#���@�I��J H�C�y)��3#nQm�}�fn�/��{( ��p^��r$$u�A*(e�  �z���o��3��@����{^E����鳪�()q+M�����cS�"�>�̭,�h�P
��|s߰t�=AJ�:<��#�}�)%� �='f��C�7#/��@�Po�I�P([���$e���$%�0��t� =�bVyqVH��y��'e&��ZՅ=dS�P�MI�Y��Ө-��ߨ�l"X�nTW����s�X�46�0�V[)��w��|��7����H��_u�O��Bb�O�d������P�2��}�4��h�I�%��*1*�g$h]`@���E2)%6�Y��+/�I��@�K����t��H�V�$���ǩ��d�9<fl$;�VJ<�{�'����${�$��p�\$ӡ�쇉?
�Y
E�Bj�+#��v��{c�j��2ɤ�K�h-ģ��l&��A5B���2��:�P,����<����hVˈ���pd��{LE�$��۲�l�e��6��7�#���&��$���H�>���[2�QH*԰�������@ h�

}٫�
B�;��үS��kcG�gP�;lt��X��
̠
�0ނ!  #�Z�.!�w8���%������did��S�:l���= F��TBXA�n�5����������30hT�h�����(���2�c��r���=��/���2�B� �%T�3�2>�9׏P}���/��[����0e���c۱:d�ɤ�KEJ�]Qe]Ds}C#���'��*�M�.Hl��!i�鋬[�5�1+�� BA˸��eDy�>���!��+%��&�utK�qL�U��V�H�SQ4���2�|;�������]�i���,��=-!�HS������J$�h��ֶV9`�dѬ�22��6H����FB���*��XYU� =
�c*4Q:+v78,3��O��փGl�)��d؏TUç�r�~��!�k���=��"�����9u6��d"_u��K��f �,{H��[��dPJ�(�� &aޠ���o{�dn�4)-.��
�Y��Ws�d|���6�r�HJ��ѷt1`1����
i;�.w7ʕ�J���Ǿ&i��^``?h�Ò��p�x$g�q�]9 ���<�*3*�dɼY��|��E���;o�� ׍!�+C�WR�|}��H	�-R�4m��(�b�o�|���d�v��w���VK(�`���A)Dq,��=9��Lp���|�u�\m���)0:���-�lv��o�����0J�C��nA,��(~`xX>۴S�0�d���)5�j�/��ξ�H��8�A�tu�N�*\n7�!Z�
�����7�e'ϓ�s�lf%]ޗ��3�^�o�97�/'���Ő��y@Zpc,1V#���������+�Ε2��.M%,0~hĸ�����f;l!����%�\bU�xvJ��1mt��� �
3o��P�4wt��sda]�-
��J���1��O�V��0�ל.J{��A�#Q[�π�=0h��n���"g̝)sk�I����:�x���oj�-�Hc[�Mr��$H-�ߍ7�hw����@S�Hk��O�%�۠kK�FCk��������D̨��T��m�����F����#�����t��fm[���Æ["��_$��Q�>�[lLi�,n���l��Ma�.��X�f0�����(] �+ʤ��T*K�RRTh��Z'��a�g$�hO���xN8����x"�PQl9���=���N���ʋ�ԛ�h#)���lS��vx`�g[�zCK���C�CxG�0@�ZC"F�Փ�v�M�z}�c-c��'���������Pg�Ήxg	���H}�Z(4�pɄN�ŝ~�u�u�YF
�x�W�Ą��Q58 �1��nq���g+8H�o�ħ��I��������9���DS.q�޹tc���/m_D�Fps������W^iG��<�E��k��L#}�9YhI�E�m�H[h0f�Z��m�)=�^��d	o��}j��U�!�(���&��`L@`8K��>�7C� �Z0�xK�n�ak�׉�2
�#�d#F+��1H+��Vm�1p`�Y
���&� ��-a����=2o����ZF��O�g�F��Uu�7Dʈ����J���6c��p� I���РF��n2�;+��E�u���
��DM(s��%��*����o�۳U�4J��1jv얂��޲�wi5�!ZL@�L0�w�y�e
���F{��=�$������.���s�F�����B���-�!�n�Arcm)F@ ��5����21ʈ(I9Fs*����v�`����R��ڦ�-qZܺ
E�T�Am���]�=����v�A5 &�-�@訊M��@�F�RC���嶥`�]�Hc`� l���q�}N�H��%�梨 y����d��5G����s�v�7��q�]�
ށn���xQ��-���X'�8!���d&ݤˡu�F\\T���`g�`�"���m�Ǩ*�7��0��܉�Ts�TB�d�(6�$��r�U	IB�%�m�G��������%�7�R��%7U�.�x���7ri�6�|9l?ՐO��3n��� D��b 0Q"e��sIm�ц7ZH>b�>a@���B6Q@k���b̝I�k≐��O2���S;�m���?�1��⫉n)HP�vn�k�/�X�º�L%J�i���p�	�'��۫1I"D��ʕ+cnH�3��f�5u��#��X�tH,�o I6ܹ\2�c�{�~W�^-�֭�Y�x�d i'7�<�8ad�1[{���(� �(��G�D�p$�	$#��P�_�B�ސ!Fs���e�5�{2F#���c3.MiG#��a���q��y��)��6#iJ��	��0��&��0��i�h�g.}�z��bef�=�R��^�6�D&����Lx��0���A�|$ ��z������]ɗM4�I0-a��^���K/ى�B.{H�D�ԟ�4�}�v�iY�p��b+��P^�KZ����y���T�x46�L�9�ׯ��)�ݱ[�:~�Ɉ�_���m���d;��}�����=�*��۶m�h^f!��[���r���������:��ۺ�/��w�o��<���:;;�� �f�V�}�RM��K�����gÆ?c�!�K�e�He�s3y72�an@wL>�)\��͹!&������ O?���/d͚5r��ڵk��q�NJ����[�韔$�(H�Q��< Fy@2��d��0��a�$�(H�Q�#' �M��S��iR|q�g���c<*I�s'1I��;��w\e���7㳑Y��    IEND�B`�PK
     ���Z�&�y`  y`  /   images/8c2f1315-cf23-4ba8-a920-becb97f13280.png�PNG

   IHDR  �  �   ��ߊ  NiCCPicc  (�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D�0գ ����d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c�%��V��h���ʢ��G`(�*x�%��(�30����s 8,�� Ě�30������n���~��@�\;b��'v$%�����)-����r�H�@=��i�F`yF'�{��Vc``����w�������w1P��y !e��?C    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD      �C�   	pHYs  %  %IR$�   tIME�WxG  �zTXtRaw profile type icc  8��S[n�0��)z^�8~$R��b;^eWݪ��HQb�0$|�>�� D�h`�dZ@�&F�Ąb�9��m��P=Eec������O8��`��Й�f�
�Q�A:���{�xt�k��7�����������-eP/���\!�����jS�u�mۃ��Qa;��B�["�,FدCl֤�	�����/�&�S�T�c��\���~�y�_���D6:J&�D�z����f5u�R�����Ye:�010�����?1:9�����{��5nH����^υZ�w�R��WU(5G�Ӫu2j�fo�-���)�:&c*+q�y&�"J��G��|/��d�c?&s&]����VG��^q���@����줁/0�   orNTϢw�  [5IDATx���w|e���3[�����!�XQ�	6�g׻��;�ӟ�SO�]�Slxީ��)6Գ��^C��m7����cӳ��؅|ޯ����y����S�y """"""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""�P �t뎇yX��s*�+��������L����>����<�r�ݵ/�ϯj>��ߌ�	�\51�;Z�w�e[�L�>��( ��R�	�NUo��W{��v��	댍
�_�f�|����Io[����7�9	s� W�>����&A����@��H��t@U���"^ n@U���^}z/[�j�[�*)9����n͚?VTV����� �*�, 4 ��{!��yLDDtX2�I�+�|���5]�dݸy����S�NMX�˯����^!"Z�SNDDDው�]8|�+LUU�S�
�n�u=&҉"""�����]bc�L������H'����ZND��fK�<�M��DDD p�ݚf���*(w��CDDD��%�$ϷX��'0���������p��a���ʓ<���#������	E��Qn������iӶ/[�lBaaAV�`�Դ48��vX�6�-fh�	�R�4J)(�L�O""":t��r�];���T�r:��'O�����z��:<7<O�����F�ۍ��*����v����"�_A��jf"��r�|��������Z�����=v�m����X5z4LZx�Ͱ�����QCrTAii)~[�+¹1k���e�E���;���^�&���� ""��:Z،m�tV��r�}^_��✕Nx�^�m�H�Q�6�5�_�6���At�z�^{�7].��#�WDDD������[u�ޤ�r9�q{"�F"""j����"b�-��t:]p{8�Q��JJK��x��.��o�\.x<,�E9�

�i*^=x@w��NDD��VPX �������}U�z<p�\�N'5C++)���r��~S�7}>*++#�F"""j� n��&"M����|��`@'""�f
�����D����>�,�E5AM	��������r��t:���(4��r� Ȉx>�N�3҉$""�������3ƌm��.�x��N%�������/ �y9�9Q���M������NDD�4 PJٍ�������(��@([�6t �z}0z������h 4��^�����(�i�ee����h�����(�iK�-W*D@�1�E=m����R�b� �Љ�����_�� t�"A��#""����+ �ϡ�ʝ��(�VZV��H�*w/D�H'����B�*�˕@LFx}>��NDD��VQY�D�Y�NDD����
��q@���;Q��*]N��!��%t�t""�h%М��J�u�h_u�8>�FDD��9�����_g/w""�h�UU���S�����G:�DDDdD��j5���~?K�DDDQK ��p�tݯCg�;Q4�b��b�W]t�)���(�i�����]��:QT�L���]ס�|
���(�i��LP�0��܉������2�fJ�r'""�j�)(���ua�;Q��bR
!:�܉���� �DD���ʝ��(�iգ�i0�OM�r'""�v͖�u]X�NDD��u*��^]B��܉����V=u��-�p`""��&uݸ�΁e������h~����*w""�����z���*w""��%���u%Ͷ���NDD�4�߯A� �+�C�)���(�i�߯��ϡE9i��5v�#""�~���J`\�.�NqDDD�N��	�)NNDD��l6[�����DDDQ�l65�`@oW�3[j^���&��Q ""#f��dX�~0�d������%سgv�؅��TTT������PJ�n�!11�������dt���D��@��!"�:��i!K�pr�V��"((,Ěu��ӏ?a�����ۊ����^�'��P�Q�4M�f��EJj*�w�#�c���5j��2a�4v":�(���fM�̡2N �ro!���b�ڵ���O���o�v�Z@��hI��� �z������ck�f,��������ӦM������b6��'�#�P\Z
�łX�#��9|Ĭ�BV�C�ϡ�I��x�d�R�=�m|�ɧض5��Q��V����TT�c�o��t����o�����_���{�]-��O7���������Wa�QG��f���x�� ��ZM�mݶ/�y�y��صk'�5�촭ܚ��-�7���Ǘ�č�wfL����/ 6j���m؀_|	�����xp�e�F:i�10�\�˄� ��n|��x�����Ͽ���"�U�&-��]��ۢ_񧫯��͛q�5� 1>�A����PXT�w�{���?�r�
��Gjj:T���d�B�*w�U����r�~�<��S((؏�L�Z���jVb��d�ɤA�4�������!�/�fK!��PX���gݏ��"�|�M蔖ƠNDQ������3�������rV�u!�a���|�8������x����sꝌ0�@n�� 33]�vEnn.�v���D���#&&�*������ �6m�m�6��
?Ȫ�ବ��g�����w/:��3�Q�Q �-[���x6oڈ��/��̀�B����F�}��nǿ��:�^�O�@�edfb�ر�:u
Ǝ���,$$$�j6n�p��(..ƪի��O�����c���5&������ks�"�S:��v8�vu"�:%�%ؿ?����p�Y X�6��҉G}���u��g��Ĥd�:}:���J�1	qq��6�|o�n�!+#Y�p�	���+0g��{�-��0�{=x���w�޸䒋�)~Y�(�(@)��ۋ �D��*wv������չs1�9�s��Q�����s�>��;	qquü����e�&3��G~�>�,r��G]{c
�Ņx���p�B��u ���B��.|l����7��ByY	�s�f2a���x��p��� !>�EA܈ ���p��31���2tx��jؼi#�{�y�UTD:눈�Q  ����]�*w���������];���t9M3��s��3�>��C��K ��f]O���z]�u�qI��g��o�e)�����.��8"�����ޚ��.@m$�q�L��Y�݋�99�3� �8�d���<1P(.*�K/����Bu"�#�D�5����EX�n^|�%���^��c�!�u�,������,7i.��bL�6-d������H��!!DBv3L�ڱK����[�0��<66�˵1l�!{LL $'&��+�D��0*�������?���9�te�:��}8��)R��ys$���~P`��f����+ ;v��']��(�O�<g�uVD��;f��8��S���/5M�����? /o+���m��������z�v���z f�6�V�f��v���G��4x?����|�=p{�����X,�Z��Y�0�L����zo��v��vCD`��`�X`�Xj�o��
��p������v�����������
Ku��6���������vC=��f��6��+_�Q�ן9p����z���`2�`�Xa�Ya�X`�~\���,=F�S�3: ������]�����f�ߚydMi��7"�^@��U�_�V�Z�S+1)_r1R����& 118k�x���QR\��H.5Kh8p� V�\�n�f��}{�b��X�n6oڄ�{������j�"..�ѣ����!''16[�>����rTVV6���dBJr2̍���/,Ě5k�d�lX��w�Fee%|>lV���е[W���#F�@�~����Т������k�d��[�{���鄈��p >>9�9:|��>�{#.6���T^Q�����u��vj����dX-���+*.����d�R�[�;w�Dee%�^o���ƢKv6r��b�0` R��[�6���k׮��ŋ�n�:�ڵ�������|��CVV6C�A߾}���|iN�M� (-+�֭[�v�Z�[�۷oGA~>\UU�z�0�͈�ۑ����]����4p z�쁄��v�ٯ��BIii��RHLH�#&&h^Wy<عs'V�\�իVa˖-�?�W�~�V�������Fnn.�����#==�6/Z���N���w�Ʉ��"��_]�QPX�������M�w8HHH`MBCR�C�r�ϡ+ e��OPU�Q�|���8��qM�Q�0t�|��(�!.>���ӷ/��!C�b�ر�r�]\R�_~]�O?�?��3�mۆ��2��kf�b��%;cǎ��iSq��ǣszzuN���:^y�U��ƛ��PA�Ν�ēO�wϞJ8�v��ǟ|�w�}�V�DaaQ��P0���ԩF�9
^x!N9eb��pj��{�|��gx�w�b�
VO��SV��;w±��/��=��9�Σw�}s^x���"���D<���Z�DFM��8����s���;X�t)
��k���43R��0b�\p��6m*R���-��������罍%K��� ��x;�iiiw�Ѹ���a' 1!�uU�G[�m���_�/���e�q����\}�j��l�Թ3����S�`ҤSЭk�6��*����#f�{����T�Z����o���hpL�UU���_���a���c�8++�)�dAJr2�)S�bƌ��ۧL��>��~̞�>��chZu�Q@iI	����$)�����nGBBB���u]�̙3q���T�� 6�M3�y)���7����DDV�Z%�{��~��i��Vy⩧#�?~]�9/�,g�s������g�Ɇ�����\��{Ӷ��p:�O>���8S��S덑�Ο��T����䤓O���������9�~�����������EV�ZU�Ϊ*y���O�-���XgBb�\vŕ�a㦠i�r{��O?�'�$�Vn'5-]���u�c��V��?�4_�R�����+���RN�<Ebbb[��������s�=_��\ix.y|>���2����kU�$&%˥�_!6mn���{��ǟ��#F��jk��^w�[m12�����?�)

DD�_�jm��x�z�.���9/6ȓ�k��5��t�Y/]-���"�ǞxR��燝��W.�����_8�9���Z<^o�cġ��������W�$&&�Đaß�L����y#�+R���_��ax�euɑ��GE���n�t��oi�t���߸Q�t�%%-�A<�">1I.��R� ~@��_��[��A�dw���V��H~a��q�ݒ�֩Z�~e�&�,�W�j��""%ee���K猬�������-r��dͺu�:���w�(ej���4��O?զ��G�̬�6c%���c�ʏ���$_*�Ny��$�k�6oGi&9a�I�h�v;�}~�|�ͷ2q�d�Z�m<v�C{L��v�Y���E��5�|s޼ꛮ���ify�ŗD�����s5zL�s�m�`���9�] �6l+�=^�\z��횏W]�'��}��|������?Q������UW�)DfBN>e�E]���b�����o����
���ߖ� �9J>��3���%��^�F��W]]�d�%��N�m;vH������n�#��n~�9���d߁�KG���Y�����n�Y���z��q�v���|)���{�%	���S&O����IgU��0�E�V�V.� ��<΁�,���x}�V�Y$t@����""��[�k���u��)S��漼f�π~hzBb��'���) ���X�|E��4�5
I���3\8�o+]�	���j����h�2�>�'PJ�j��j�C�����߭²%���k����~��#L{�R
%�������˯�����뽤�>5�9�K�����|�p&�y��g�tVɳ�o磏>ċ/�����������O<�gf?ge�i�k�O_Kҫ���O=�J�n��=�O<��#(+-#���?�v���k<��l���V���³�<�[n�۷�ե�����Vs�����f��>��Ar���5����Ǜo��nǲ�O?���|vl�Z�/�Ϥ���`�5T�����<���t����ԍe�7z�����c��
�Z.ս�Us1��d^}���طo���v���T����	۟17�p#�6oBM�4���cࠁ9r��� %%�����{����e˰r�J�߿��3X�sN��my����a��q�駵S/V�߇���:�x����n>�c��ХK6z��.�]�*W�����u�VT��:F*�~/��70}�t�\�
�̞�*���vLGl<r��W�^HOOG||<\.v�؉u��a���՝Ϥ�qW������8���o{GB����x�w�rU6�?&�YY��ݻr�� !!n�شi�l1�	@M�2����8��3P\\�G~�����=Ɓ��������HLH�����]��~�z�ܱ>��4źߋyo��̙31n�Q-��χ�^~�f݇Ғ"��:�q�ӧ/F��A�!5-q��p�\(,,D^^.\�u�֡���^fԧa��������O?��G�^�+��+V��9/4� p��!;�z�쉴�t$&&����@����!o�����=�7?�}�]L�>S&�2=�z���Q��i��z�oټ~_��ٌ�}� !>�i�8�ѣG�ꎀTK <d�ˡ�ܭ�yu�kQW�|�_""��J�R�� ��]��E�qy#"�l�
>rt3U=��N��?]#��^�
���Kc~]���b��_�o7��dee7S=	�?`����/-�[�*wM�[u�w���b���㏑'gϖ�+WIqI��=��|��z���R6m�,�ϙ#Æ�Y�e2Yd��iҳw�F���O��N?S�xk�lشY�+*l���T/]&��q���t�?&�U~��v�r�+P��0_Lf��5Z|�Y�t�KU��V�\��m�����2n�1�4S��*M�Lr�Ie����|Qu�㈓I������%kׯ�����RZ^.+V��Y�= �z�}�(��|�m���Z|ο�����_�?q����k�u��r�%��'���?�DN;��z�����������q��R&INN���uHjZ'9��d������������|�t�d�Ν��G˹�/�	I�^�:�).-5L�_MP����{���={e���7ߒ��� �TIrr�����o���g�����҈_'U��_­rOHZ��C��2�[��ʫs����楗_��fx"6\v��uD午HQq��w��m<�����O?�J���bj�""UOu��)�e����8M���v��
����j����Y��n�^�{<�>Էd�r9���͗���ӷ����\)*.iv;^�O���2h�Аy3ᤓ���(�1
���%1)E���FٴeK���˺d��[��$�kwyj�3�?���|��|���d̸�C�ˈQ�e���a狈���;��ԴN��{�!���m�\�����By��g�i�V2��0��)bЛSM4�E�?a�|��gRVQ��^RV&/��buڍ:�)霑)?���;��_~)���Azjj�|���I(��VFe@4x����^y��d`mF����;���I��������W_{Mb�/�J3ɔi�ʪ�k[��""�����s����Dd�G{\���N��E(K^z�U��x������V��s�ꐡ�F�7�~>��|�駒��E�j��v�!�W�{��z]�$����O>U{�nz��Xz����Ss���ǟ��脻��� =z�6؎�������~{��*�\w��B��Kv��2�5qU��[r�麼�����|�8y�ŗZ�
��,\��?ʖ�[�F���뺼��[ҩ�q����Ly��k�9�u>~u������8�����C-�˴��T]�;ŉ�����:nt��	�6�m��{�⥗^FeE�&��0�$<���n� �z����>���f���
��}6nl�����o���a�X��p���>}zXKgfu�=��N8����:e�D�v�ü)(����[�-W �l�⪫��UW���E�2b�p�}��P���>�)�����1c���Z0@� 8��8�����PRR�6��>�ſ�ݷ߁H��i�Ĥ�~���a�Z[tk�z1)�3�8<� :gd��5E���ܹs�s׮��Li�y�L�ݤQ�^����:�L\r�%PZ�c�������QYY����tPi����,p�W����LJr2,Cf����,]�zZ������v+���ݦ�5;��~+����k׮Ň~�E('�|.��RX�ՊI�&!>>�B���p�e�a�)���ՊSN����S�*T���eK{tcǍ��W�16[���I�p�ĉHMKCs=��=�\�}��V.��a�ē���t;^��7o�?���U�|�-�޽��wM3���/�%_sn<�	�g�v���
��֠��t�̟�em�ӑ��7�x:��55�%i�Z,8��sеk�n�桰��]RM��iF�]�H������^�Fb�#��eYE>��C��A߷Xm�����;���_#G��u�]�#�.c�ߋO>����k��� .>]t�SS[�@VV�/�:�v놙3ς�ln�vrs�"-=x��u?���ۜ#5�b����.@���V��O�>�޽[�|t��s�;���k �ٳ'��2�#(..��o�͛7�/�2X�����_	GLL���V��^z	�`�tw��~�	J��ڥ��4Κ9�n�q�>}0d�P��K��Q^V����@4MӚ-��,�+ >�����餶�>o޼K/1XBG߾}q�9g7���-���N��#G���5�VW����_�~?��6�%=-�YY!�9���ѿ�6m'%9ii��RQQVI4�|�ޣ;&L8�MkINJBN׮!�3f���)�@bB:w�l�LEE�z�!�����m��tn2Yp���!77�ݚ�@�=0��i�M���8�&��֩SgL�2fMk�Ͱ �����`�[e����+���n�t́et�������v�M�h�"�ݻ���5�<q"zT�õ�ѹ3N�~�aUdYY~���v	^�G�F�N��Plv;:g�يѣG���>�ݎ��$�������|�0�aÆ!��s`�X���a���0rԨ�Y�ZC!0�_rrJ�|q���1�� 2?��#��`������ĉk�@m/&MÄ	�����7������Ö�����>�+jJ�k׮0����|>����5���DS��b��9}��d��zz�`D�6�Jm�>�-[fp�$��`ʔɭjwn�0q����%���t,Y�eeem*i��V4���`2�[=�i��JHH@�v���b� 6�a����m��3�L8hP��6[B�4����h�a�Á�i�@����.��y�73���}��r�*���>}z�)�F��h���<X��o��xڼ�A�!11��n�SRS`���	H?����%���xU��HE�{ȥ������
@iY6n�h��]�tA�~�Z�w��}���m�6��o�1z����j�����$''#�Kv۷c���tٶ2��j��w�^mi�v�a����ѭ[ז��`;m팚��{��Q�����Ў��� �d�\ߴiS�o^�2�W�ۯ1..��fXD���F��@��r�4MCL��4�i��RXX��;w�߳WO����l����ܾF���cZ;w�j�V���;����iƗ۸��fn��N��:m�v:��m�-�)���X8���(_��~õ%/�e���f�w�.��c��{�n0��ٻg/���߆���vdfd�9��X���ۤ@��TbVJi!�H��J)$��#T�����6�5�G�����W��Ē����؃�̽�d�`2Yj'f���҉��m�F|\<�����q8���9 �)�@�MHH8��c�=D3V������m[�3���Lطw��vA�� JKK���ڪPR\��6m�j�"9%�]�n6��B��v�8m��T�w��)�.���Lf�����t�x��hTPPgee��Lf3����Ih�tɂ�b����$
~���-�;b�i�bs����j|��������l�Z�'���<��~ط��MK�^�O<�8fϞ��-Q�݆�U�ۍ�¶t����G����6��A%f���n ''6�.��N���p:�H	��pQVVVݩ��~
L��z ����d[Uմ)C�u������j6[`1�@��:%��c2���RZ��mP <^o�APD�(5M����P\ܶAZ4�`��5��2�B���9�+ ddd">DUdQQ
�x'-�n�a�f2��#�Q݋�)A��m�Ř�&�ڱ�Б�d2�|�^�V^OscL ����+8]U����J)��C7k��nGm��f�~�m� ������xRTT���o�]�K�1w�*@����]v����9�`>��M碦��E�p�iLGؘ
���>x=��E�"At�vxl�:i��;�q��;���O߾�FGZ�fmTݙn����+QT\]��(Tk���_�W����Y��Pe{�T�����zЎ���@�����G��e�h~������.���?�Ƞ���ʕ+�t���=�����SO>�?���r1l�0�9@NN`2��f����_�QYQ����r��	>8��4�cbjg�"j��M���x���;�<s�O6�f2�K�.�%:�����r��G:��� �>qqq�(����+�}�h���ښ�����_�k�v�ڵ�|���t��@��}0b��u֙8jԨ&�)���i@��������"�t�������QS�z���1��!+���s_������f�s�7� $�znC���#'�+֭]��]Î۱h�t X�~=���P����ʅ���}[�[���郣F�j�ل��m6Tx=h�Ș�������������mSi�Z?8P=�Պ�x�N�U.bc�پ��&�D-��U�!���`����wW�������rE�u֯��n�w().F「�1�2220|����OMI5|F���b���}�m;vT�����l6dtj��̨c3��HO7��N���E����$�/��f[:n@ v��'MBl\��f�-X�e˗G,�
��m��駟AĨ3�`��a�ݫW�w�;�W�����P�t���ׇ���A׃����S�N=/��g�n�6S���;w�t2�ZLucu,��ƌ9
��r��$�iؽk7��{��ko��9֭]���M�7[l�x�)HLH�SSS��c<�Hޖ-(*j�`F�Ôb��͆�$%%��8�D�޽z�f��������o���\�լ1��҉�&��Ն�1�_��.]0i�$(ͨ׫�?��.\tȿ�
���7�xOU]���G�8���1!!}g�Rؽk76���v۶m���[`ti�ѣRSSbNRGҳW/���� ��%%%��}�Y_޶mX�b�nۆ��b������ܩMj&
���a�4�}�L������ְs�v<��c؟�Ⱦ�
�����9/b�0�7�0u�T���ǰm�j6c��Q�XlA�TTT�/�����m��W_c�޽~:j>b���ٶH�{�n�e8߹���k�j��v�n�Tŷ�z�N��3N�g���/�7��x��G�漷QTT��N-"�hh�U�w�*w0h�@�y֙P���_|�^xa\n�!�2~��Wx��W��U������9g�k3�{�1�32��E�W_}��۶��) �������/t�}���aԨ����$
� HMI��1c�&X�����7o�m�/���|�}{�`������x��yx��'q��7�GCE���!Ҵc�:v��b"�Й���z���O���SO>��^zn���u���q���`�>��- e�̙ga��ͮ�o�>}�h�w5l\���|�8� ���ϰl�2�}���aÆ�ܤ�Ƥi8�	HI1�Y�g�~�%K����X��t����7
���!��W`KcƎAff��L&4��XE�9�zˉ&�t�:�s�u�(�_����fw x9�������栢��u��E���K/��=�����/���)^@B\�O�{L�q�=�*<������e����Vᩧ�Fee��{�2aڴi���>�/pth�5
�F�B���a�x��Ǳw��6������W_ᓏ?6\2>!	'Nl�6�H��Ï��5d��i�pJ�S �Ʉ�.��N��C��� ?���|˭؜��n]m�n���G��O�`ѯ��X� 6.��_0hР���ĉ'W_��ض5�� �mk�>) ���C=�իV!xէ��ݻaƌ�T��UM��y�Gl�:�}��'x�٨t�~������u������� F�Q����C�{q$�ڬ0�-���'����9�L��@zj*n����ۯ?�= �P^V���'.��b�2�5�;�ߪ�^���<�}�?p�����K~�6�L8��p޹���, ���p饗��Y澜?7�p#6l�ܪ���k��r�mx��wO0�ɂ/�C�a��iӦ�㏇ѹ��z�ܳ����BQ+{�+z��q�X��Q�UABb2.��rtJK��{�#6[�!x<-Z���΁-��7�_¶�z�����u'2�d�8�+躎_�	�^s-.�݅x~΋X�n=���-�����+1��q��s��#�"����8�N��[n����P�8�t̘1��}]��>�5�_/X �����Ѷj������E���ÿ_��M����
Ǝ�+.�V���$ux�SZ���/��2�.+����ч�M7݌�k�A�0�58�u]���~ß��>��Ð���S&c�ē#�-�L\|b�1�
�}�̛7e�+~]���g���>_�8?3�M)�}��pV:q�m�#��>�zd��t⛯��?���ݻ㨣�°�Cѯ_dee������NTVVb��}X�b%�/[��K�b��mգ�5׏Q0v�8<���գG��� HIN7ހ�k�b�eA�MAD��W_a��u8��p�93�۷/����҉-y[�чa�k�a떼�u5��[�����н{�QZ�șp≸��k0��Y�r9���T��rᕗ_������/�ӦMC�n]g0\���
y[����c�ܹؼqS��<t����IhR������aÆ`�*�ٳ��z����0` ���PU�B~~�?����Zx�_C 1�|�fo6}>�9��!��_|�Ep{<���b��=]j���x�i�zlڸo�a���@bR�6t�\.8�NT�������P�a��`�1������#Z}����1�Y����my0z�g��]x��G��o`���}�hdee!55&MCaQ��ۇ�K�b���عc'�~o�}ё��	����4q�8�ԁ	 �ł���
�v��K/�T�hӠ.��5�W��nǜ9s0|�p�1�3����Ʉ��r�ܹ+W��o�-�֭���y�|�;�#G�0�Y��=z��g�T���G���>� Ji���ǟp".���%%u�<�����}3j�\���
t��	��+VT�*�_l]�QQQ���2��j*��i�-VL;�T�{�=<p`���S�L���p�-�`[�u���;�g�N|�駰X,�X-PJ�������DGVv�����.�I��e��N �$%���^��z�MA�^/�lڈ-�6��wޅ�j��b�����v�ü��93w�uN�1#�W&ҙq��l;v,�5>�a�� O[ri��(,,DrRR�w#z����yUs����eO� j��̳��+�����<�����	��^��=	w������sϴ[0 M�0s�Y�={6F��y>�h�u.��ge%*+*��x�*ԅ-��!C��SO��/�����ړ �����܇��+���{\s><n*+*QYQ��*Wu�i�|��={��G��W\���!��I�N��aC�5 
�����H'?�h��;����Ç���O>�����b�"p��|\�q�2�T���+���;�����[Ӕ©S���W_��.��	�a�W��*���HLJ�e�_��_g�y&,&Z��[�P�+�j:��}�]x��'0t�(MC�`��@5�K�|���<�T�y�E��y��ͭ;އ��.L�s󭷠KvW�$�WTT`ǎ�ޅhn:zs@��4�����)���{������5kQ\T���Z�խ���̒�����1c������ɓjs9XGH <�<3�'O�+���E�����%ψ��GRr
�=�X\tх�4i��ڶ�n<�t�i��� ����4���vj�_�01�N��K]�������X�����¬�z��rI��o�V@lL.��b�;��}|��6o����=?Z�y��5�����_r1.��|dt�Ԧ�]D�=��ů��~=	<�l{��ߪ���f̀���+W���>_+ۨ�ra˖�����ݙux]g@oV�i�='���:\x��X�r%���{���ö��P\T��e0�w0
���I�ջƍ;�L:�F�DjJ2���
s�p��c�ē��w���>ǢE�k�.8t�N�̈��C�^�0��q�2e
�9f<��{���S
�9�2tX�1�u���ܾ0�ZYj����l2��HW�_G��}`j�H_�@�G��1x�Ph����޽{u	�y�6|x�s]ב��[��v���:lx��뺎~���j��b��(���9��_�ѫWO�Z]�S�f@n.f��\x���������`��U(�/���Fs%Jbbc��)Ç����N�	'��ݻäT����d6UUU. "���T8z�V||���Ғ��/8b㐐�ت�6�L�y֙0` ޚ����%��塬��6�( J�`�48bc�������sЩ:�2��w�ݳ;+��_r)^x�y�m6��@M��"(,,Į]��c�l޼�7oF~~>�N'\�@�v��M�`�ِ��Դ4dgg#77����ӻR��`�>�#u,j����Ǝ;�n�:�^�[�n���P^V��
����@\\,233�77���b�����̄�:��~�ʊ
8�Π�[,$&%Ak�ޝ��p��o�j�"!!�p���G���vv����\�W�t���"�{f�III��p�Dee%*&1�-HJJl�픗���r}/��I+_�Q����Rlٲ�ׯ�ڵ�k׮�w��n���!6.q��HLLD�޽1`�@���=�wG|\��;߫�n����=�4�II�߱���xQVVt\�a����M!P�p�@>��m�Ν�p����N@)���!11	����YY����n{}D�_�7<�ԓh�&4&&f����ڳo���P���]��^z1v;z+��]A���x<�z��z���|��|Д����
{LlVk��F��g���������J�l6�b�"�no�6~����/w{m�p����hَ�6u ^�.�^�70��R�X,�Z��Z�������<8X�>(��ߏd-�fa�! ��o�4���p���~���9�4>#�&���b�u����3�Ѳ�m* V�VKBȠ}0��<8�ېF?��z���ЯlCoo��k?�N^�)ԑ�|?��kᡦ��|	��:Q4-�����p�""��$ 4�ërg	���(J�Hӧ2�E9	���e�8""�(&�.͏3�6t""�������Q4-�����:�E�:�5_B�u�����(-�)�D�˝���;���0¿�h�DDD�>�.��V��0�E%DCm�::QTif��z2�E-�$�6tv�#""�Zv/wщ���VJ��DDDQIDD����Љ����ha������(���;#:Q4����3�E)��{�����(j�7�+{�E��&g�s�DDD�K­rg	���(��`�5��E��̶�Q0"��Љ��� ����ֈ���Z�Я�U���;Q��yl��`�XNDD�D��|l���(���Y�NDD�D���NDDtؓ�Oe('""�ja��V�E�0��Y�NDD���ǡ_����[���8�+Q���H�����Ba�;��#�8Rё ���,�E�p��YB'""�b��rg	����c,�j-X�����Vؽ�Չ���V���Y�NDD�X�NDDt`Fu""��ő∈���2s""�(��ʝ����NqDDD�?ζFDDt�p,w""�#B�m��DDD�,��eX�NDD�Z0�E+�GDDt��ќ��(J���;�Љ���Xx%t�r""��֒��։���T�c�3�E%�!"":"�߆.�r'""�V�V�3�E��*�棵��E��c��Z�)�����Yx%t�C'""�R�oF��Z5�ADDD�R-��>s8K�u���()-�����C�D:J!���h]ס (��4�]���������*�]�+@s�	���jE������U�HD�Q�y����>x<(M�b��d6!PFm�밴�����ػ{ws�U���J ��W�1J�DDD�C!�[�* W�߆v�'""�B���Eo""�Ù���G:%DDD�j���tJ�����t@y5�ie�N	�� ���v��H�����ZGӴ����2-%%�q�Ų������#�aK)����φ��F@Ff�q���wy<�" ���j�U�{N�p0:�%@��iͶ�����pD�g?��������9ETM)��R�V��}gm\�a�:����F�~�w��ի��2"V f��b���1&�ɪ�4��4��4�R�T��`B৪��R5WE�T��k�U�f�.�PX�v����RhxW����x9.����R�<\(T�]�R��ԀR����u�V���o5�k���^�=�:Z���Y�~Ԧ���������j��d}J��u�������4��Z��p�	��ʂޠ��^��u��c�o�5��b�x��/=��WD�H�����9��:{�~���������nHBi�{ͪ��R�4����k?���F��w���'��f�!��`geI��5�|M^�~�������4�	��t�cP��V�p��Vw\��n�f�'�z}���`����~i�'|�P������e��e��FK׻�68�W� ۯ9$���dݵ��p����u?t����������K�Y_��]�j�GR/���\�dX �5ikt\��*e�R�p��I�ɋz���ͯ?��ڹ};�~x�W��]��E��O�����FGT},�4��o
 �t]����߯ ݯ+]~�_��D �_W��t%"�~��s��oP՗]��^W�i� ՜ "�7H"XMŊ��>���]���>k��כ����}{��m�9��g���_y�7���4������]�78�J)���x���q�I'��^O���_��5oIݽj��O ��V��b��Ҡ���"5�RR�����R��$5W��;_���U_���BW_]�҅�r��ȁ?���M��r��7�R����d����/U�=}��Li��i
J��MдڿiJA�(/nKE�c}+M� Д��Ai�mk�Mi  ���;�ݨ�j�,��Q{JNIE~�<�쫇q1� ��)[�fʼ^�}>8u14��4��~�AY4(� ~?4ѠC�I5z�_�h�P ���\����k�R
���5��=�j���5�^[k�ª��5�)S��/uWߠ�cG��ɧLz������-���+��s�|6��0٘PRZ��n�/��r�������#F�87--}魷��ߏ�1���d�l����&��-W�ƥd�hT�Qu�T����7��n+�ꭣ�i�h=5�u ́�Oլ\I��������R��ڂQuU��K����[����_�D�N�	�ʹ�p`E���Hmy]�4����P��nOS
�i]��L�u@��lF �X`����*������t�	�v#..J)j|����Kv6X/�y	&�����D|B��v�G�7p9�� Æ��m;v���."�Ꟈ�����?"1�Xi����*���?�㳟�[��E�05�ک���L8�$�������M�Pغu֮] Hk�a꣏?�?���`��������'���Y看��6�sύtr����w��w��[o뒙���a���Lr�=�8"J�""�,\$	tMh��q�ۏ=q¸�YY�>,DD�XB��23�0c�i11��A?.\��Ҳút� l۱w�u֬^��_	������~�o����[o�S�<�$ŀNA���`��1n�ñ�d2]f͚�ض}[���j
@IY|�!|��Wh�p�RSS�>��c^�~��k�N\w�5�N6Q����[t꜉�cƞc�����ݭ�ye��ڎq������#�=.��xi��O�ظ���=�8�#.҇���Y,�SP����٫���7[,֢`�x�.��˯p{�	�>��3<��cpV��q��d6{323������7�Ήtr��Bb@���:�����:u�e�Z����l�2���V��
��U�qｳ�o�n4�(�����G5�I���6nğ��C��MDD�:�>����k猬7��t����N���?6��""���Η���ILL���#G���8"}���ڮ� ��={�]��A���d�'��}��*�G�w��l1A��M&�;;��"���.�sϽ�>DDaa�;��q���d6W[���b��%�r��j�O?��>�,�n����aC_7�Xٳg���H'��(,�d���>Đ��Щs�-��Ш}���8����T�n~߬�p`�^;��11�srr������G�?yB��MDD�>f�s..�������_�UQJRR���oDm���ȁ����f��٭[ϫ����/��F�����EXB��F�����,��>0�}c
%%%X�|y��j�������G|�}�)$%'�w������S&cǎ���D:�DDD�G����?`Ѝ&�E^�����rE])]D��>�N�A�i4��KX5���t���&"":8���[d�tØqGO���F}��a�u���	���`�|�J>r�a0�X�e}r�] ��}���NpDDt�:u��8�̳�&$&m1z=)9U��u������!�͕f����go����s��_o�!�YMD�jlC�f%�$#77woLL���K(���bٲe�Njuj �׋�_��?�F���0��~�j���x��"�t""���G���={?��I����9�|�p:#^Jy��s�vs��Q0hȰ �~c,X�l&"":�j:�6��f��g�"[�n�h@�����#Gs��������w?��r���]wϊt|_|���O�p��Wh�<zbb������v��ϛ����u�ge�?�x�4qR������й�Kq�Eg''��
�5Q�$�=�`Ăys���8�v�=�x(3���"�Ý9�	��CRb"����6
���˖.���D�ÁC*?��x���vW!�8�f�ٓ�����E��p�ݳP�*�R���DD�c/w
Kf�,\q٥����U�f|ڬ]���8�iS V�]������A�`��BrJ��G;��S�L����x��q.E�� �KF�;�j����GOLJ���y���ED
���/(�v󸸄���3<�s& ��>�t�z_|�N�p��:}P|B��P��<��#�$���x�^y��G�k�nn������� j6Q#�#��),�'O�裎����8�-'�K�.���:$����xꩧQ�D��vMӐ����i�Ϙw���`���8��#��DDD�ܜ� "Z�^}�`f�a������^3N���e���>o�IbRʢ�&��k��!����,$":hXB����J���V��f=�R
�v�Ė͛Z:4 %eex��G��/���4���]�u���W_nY�|n��o��B""���>j,N�xʉ�ظ�6kM3�#�=~�J�^�_�|z�8b���M&��[���������\�;�~O������s����GϞ���o����묬L��^ݎB��ޮϣ+ �}�=�x�	8+��txD��Qc�z殿�����>�L�����(z<�������]�u��xxUȰ�#dێ�ZJ�ۺUN8�$�vsh��m��㏱�c  o��v�����(��߸ 0pА�4�,Fϣ����7�k��."RVQ!�\�g1ޮ&��շ_������{���#�eDD�;�Q��ر		IHNN^n�Z���R(--��+�m�~��ƛ�׿^����oUӐ�)��S&M�{�Y3e�M����t�E��3N�̳�����ۨS ��K�UU��R���?�$��䆬jOLJYq�)����,"":�XB���������p�n�ܚ�kPPXئm) ;w��}�fa�0|D�n/�޽�_9͇}�����HgQt{� "澹�_2`FIZz'��ZUB�W��t����ILf�a�\3Y�n�{>�ҫsmW��Z<=��HgQ��UU �3�:�ŦZ��*��}��U�~y��Krr�W�k�����3g��3���0y�4�qNDD����
#G�i�Θ�P���+/UO�K�""�M�����=c�>�d �DDD-u�5��ڿ\ףS�����Qc�ɞ���.�׌Ӿg�>�q�!K��͓�o�-"��v�x���"�-DD�Nq�*��;��O��!�U۾}�n��z�*��>�>����S
��>�0�9g�9S߱s'�v�u��""���[�[3���&�%T)Z��R����󎤥wY:OLJ�8q�Q�9�  �/�t�~D=z���i��pĹC{՟�������V����G�l7����G��= |2�K����HgQ�qrj�-[�`��G#..n���(v:+;U��^���%蜞f8Q��_X��+�-�Qk��i�ҥ�[����7F��5�V�9-*Q�=��l�~{���[��qY]rdђ%!����̺���cBV�wꜱ����;�����@���������7ބ��G�>�ߡ&j��b���n�ED>������jW���P|܉���7��>�t����{ ��S��d�;ĸ]�u��M�>_�`�f�:9j̸����M<t�c?.��z�?f��g8�9Q��vƙ��UW����^���ēN�����t�������J偗R&�ֽ���xc��睏��^�]'"":r�����Y���G��ޣ׶P=�kwY�|E�������ǟ�G\�vs%)�i�Κy�$ p�uk�ϵQ��v~[�,��1�~0�r��~�?�Ou����_~%9]���jWb���{�	w��魷����|�]&"":򔔕AD���N�b��hG�t��]���{ٴe�{�	!{�k&�<􋧞y���7܈y$һKDDtd��変�\i��xC��%3N?CV�['��j1�X6;���k�������W����G��Y����}��l��\@��8d����h��<!1�s����$"�_~����#��DDDG�5k� �Sgddgǚ��OB�������Ymr�	'~4��S�}�y�:�_��M""�#ߥ� ���z�����u�׀���=����:�\ �眈��8q�46�;>#>!��s%�]���DD��nl޶-һGDD�q|�� ���g���[��f�L�>��=���~��7X�zu�w����c���7��~������̬�ו2�8��cbw�vƙ�fv���v""�����G{܈ظ��-
�J�9b���õ֦�:>�/һBDD�1=?w.�="��=z]g2[��	��"i靾0hp����b��a��""��������N8��8-)!1�悹R&;n�޻��Ǥc�;"ªv""�H[�`  ����{7[�뫫ԃt�-��w]|��h�N'�{��H���o��S�L �쎋�L%]w8�^�<uZ����GT:��N:���@$%�"%5�j����i�FU��j?5�Sv�,t��k6l�t�����1�dA�Ι8pprFf������Ė����LIM�ӳOߞv� p��wG:�DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDG���Nþ�C   xeXIfMM *                  J       R(       �i       Z       �      �    �      o�           ����   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��    IEND�B`�PK
     ���Z�����  �  /   images/6fc4b800-efc3-4a5d-827d-9566cfd108b3.png�PNG

   IHDR   d   d   p�T   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK
     ���Z
�8b  8b  /   images/a7e3301e-fb46-458d-916f-a05c0bde95f4.png�PNG

   IHDR  �  �   ��O3   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���]l��}����%R�(��(�"mY�-?(˃���S�$]Ңht�:l��u����C�m�i˴�Л]�z�a7	$C
�hs5�r��b9�]�ReZ�����"��8�BQ<�����z��s>�o��/S  �laa�G�"⹈8Px� ����N�*=Z�7�7�^(=   ��.Eę��}��� "6K ��T�  ���=�"�E�gC�     t�LD|:���^8z��J ��� xU�s���C      �ӓ9�?>z��ϖ  M� ��������K�      �!�9��>??���C  `��  <P>�R���w      찱�����=Uz  �� �I�."z��      �TUU���8Qz  �� ��ѣG�^D�.�     `�����ߔ  �"p �����8�s���w      4�_=z���G  �0� x �u��#��;      ��9/�  � p �A�"⟖     РO�����  �iw  :onn�q��     �&���Xz  �4�;  ��R�g�7      𩹹��,=  v�� �N;r��#)�ϖ�     PBUU���  �Iw  :������     Fק���*=  v� �NK)���      JJ)���  `�� 謥����;      JJ)�Å��=�w  �N� �Yu]���      Z�@���K�  �� p ��r���     �6H)���  `'� 褣G�.F��K�      h��.--�(=  �� �N�9��     �6?_z  �/�;  ��s�L�      -��  ��� �E���'K�      h�g���N�  �C� @�,,,<ӥw      ��`0���  �~� �ϔ      �R�Pz   ��;  ]���      Z�������#  `��  tʣ�>�;"�)�     ��R]�~.  �%p �Snܸ�LD���     �bw  :K� @�|��      ������  �!p �k�      wwpaa�åG  �v� ���     ��L�  �w  :c~~���8\z     @��?[z  l�� ��H)=Wz     @���9v�؁�;  �^	� �ӥ      tD������#  �^	� ��;     ��?^z  �+�;  ]ы��Rz     @�|��   �W��  `+���zO�[UUU���݆Q��������p'ccc�k׮�3    �j}}��az�ȑ#�o�����C  `�7  tB]ק�z�~����1111>>����v�~����cccQUU�z=A;���<fggKπV���?O>�d�    [���q�֭�y�f���ō7�ڵkq�ڵ�~�z\�v-rΥ�ދ�~��\D|��  �*  ]�����XLOO���t�߿?���SSS�gOg�     ;dll,���bϞ=q���;>���o��V���ƛo��.]�˗/G]��ݺ���C� @�� ���LLL���|������LLMM��.     `D���8t�P:t�����|�r\�x1.]�/^��7o\�#>Qz   ��;  ]PE�������Ǐ�������     �]�^/>�~�sׯ_�.�믿���zlll\��7B�%G  �V	� h����G��ޭ>_UU;v,�񘙙�4     �199'N��'ND]ױ�����Z���q�����,..>�ꫯ�m�� `;�  ��`08���RJq�ĉ8u�T�ݻ�     `h����������ӧOǕ+W��^�������J#��pD� ��;  ��Rz_����8p �}����      m355SSS��OƵk��ܹs���/�[o�5���9�DD�ǡ�  � �;  ��s~�n__ZZ��~������     莽{�ƩS��ԩSq���x饗��_����}��҇w� `���  `��^_8~�x|���     �6==�>�l|��}�C199��/�����=;��  0,w  Z����c�؝�v�Сx��g#���*     ��ؽ{w<��S��}.>�āv�e����x!  6g. h�7�x㉈�u���>}:z�^Ë      ����8~�x?~<^y�8s�L\�zuۯ�s���x~� �p� h�������gggcvv��9      �{��cii)���ę3gb}}��_#���� ��� �vO��sssM�      (���x�������g�Ɵ�ٟE��^^���  ;�*=   ~�������ɦw      �{��x�gⓟ�dLLL��o=y�ر�a� ��"p ��N�      �6�����?��1;;���ҿu�����  ;A� @���x�N_�r�J�S      �eϞ=�O}*�����|J��C�  �M� @k-...Dľ;}mee��5      �������x���o�q�;  �'p ��r�'��k/^����&�      �RUU�},&''����  t�� �6{��="��_lj     @��޽;������9��GDjf  l�� �6�k�~�ܹXYYij     @�;v,�����ȁ������  �!p ���q<��󱶶��     �V��*:t�gRJw?�  �	� h����������矏����     �j9���SM�  ��� �VUD<������<������-     �k0ĥK���L��Ɇ�  ���K  �;YXXX���[}��W^����|�#����5     �����o����]�I)�� @��� @+UUu�^�+��_���bmmm�      Z���_�o~�[y��� �b�Y ��꺾��="bee%���/����NO     h��^z)����G]�[y|����C��  �%p ��rΏl��޸q#��կ�ٳg���      �s�ʕ��?����7�qO'�����,  �/��  �NRJۺ�~[]���o~3Ο?�=�\LOO��4     ���_���ַ⥗^�ֱ������/��2  �w  ����._�_��W�G�~��111�/     Ш�s\�p!�����������>�S�  `�	� h�	�#������w������O�O<�w�ީ�     �����p�B���k�ꫯ����N��� ��� �:���;��q�������'O���'O��     ����f\�|9.^�.\�����x����  ��  �N��{h�����/��b|�[ߊ�z(N�<��[     ����㭷ފ���������t�R\�|9�n������YYYy��7 �{!p �u��Zl�}꺎s��Źs�b߾}q�ĉ8v�X�ݻ���     F���f\�v-�^�������o��V\�r��������c!p �u�  ��R�ox���8s�L�9s&<KKK�����R�s     ��X[[��7o�͛7�ƍq��ոv�Z\�~=�]�kkk�'���"���  �&p �����^�|��x��7�^�]�v���\������L8p �}�F    �����X__�[�n��������vȾ��7n܈����W��GJ��  �N�9  �Q��������{��^|�{ߋ����bjj*���SSS�o߾����ݻw���x���^     �����9G�9666""b0�����u]���f�����ǃ� ����3d���,�?�Qu]� h%�;  m�Tz�{��:VWWcuu�=���z���\���c����X��J_��W��ٳ�g    r;Dg�\p ���  �Qk.�o���/�hx�(��ݾ~   @+=)"r�!  �NU�  p���     ���\\\\(=  �M� @����싈��;      F�c�  ��	� h�~��z;     @��� ��� �*UU-��      0
RJ���   �&p �m\p     h�#�  ��	� h�;     @3�  ��� ��Y,=      `D/=   �M� @��     �1}�����G  �;	� h���      Fŭ[����   �$p �m\p     hH����  ���  ����̾��*�     `T���  ��� �������      0J\p �m�  �FJi��     �s��   x'�;  ��RZ*�     `ĸ� @�� h���      F̱�H�G  �mw  �d��      ����ѣӥG  �mw  Z#�t��     ��Tz   �&p �5rγ�7      ����  �6�;  m�;     @��  ��� �6�     4��룥7  �mw  Z�رc�1Uz     ��I)�� @k� h������      F�� ��� �
u])�     `D-�   �	� h�^��;     @.� �w  Z!��;     @�=����#   B� @{��     PH]׮� �
w  Z!�,p     (dssS� @+� h��ґ�      FUJI� @+� h�     
� �w  ��w     �r�  ��� ��p�     ��;  � p ���8Tz     �� �
w  �;r��LD�K�      aK�  @�� �v�-=      `�훞��*=  �  ������      0�v�ڵXz  � (.��;     @aUU	� (N� @q9g�     �[*=   �  WU��      �� @qw  ��9.�     �8Zz   � h�;     @y�  �� �6�.=      `��gKo   �;  m p     (,�t��  � �w     ��\p �8�;  mp��       bbfff_�  �6�;  E9rd2"�K�       b||�H�  �6�;  E�z���      ����gKo  `�	� (*�$p     h����  %p �4�;     @KTU%p �(�;  E�u-p     h���l�  �6�;  E����      ���  %p �4�     Z"�|��  F�� ��\p     h����  %p �����      ��;  E	� (��k�;     @{�� @Qw  �r�     �U<�裻K�  `t	� (M�     ���͛�K�  `t	� (M�     �"9���  ]w  J�     �H]�GJo  `t	� (�駟�{K�      �/�z=� (F� @1+++��     �L��w  �� PL���     ���  #p �����      -�Rr� �b�  �$p     h����  #p �����     �}\p ��;  %	�     ��w  �� PL��@�      ����H�G  0��  �R�*�     �16==���  F�� �br�w     �;Tz  �I� @1.�     �SUUӥ7  0��  �s�_z      ?*�$p ��;  ��]p     h'�;  E� (&�$p     h!� (E� @Iw     �v� P�� ���      -T׵� �"�  �ҋ���#      �Q)%�;  E� (�رc�""��     �	� (B� @�n��_z      �I� @w  ���zS�7      ��  !p �����      �%p ��;  E�     Z�PD��#  =w  ���J�     �^c333{K�  `�� ("�,p     h������  =w  �p�     ��RJw  'p ��     �M� @	w  �H)	�     �M� @��  �;     @��u-p �qw  ��     �ޡ�  =w  �H)	�     Z,�t��  F�� �R��      �]M�  ��� P��      �&p �qw  J�     ��� ��	� (E�     �b)%�;  �� PB{K�      ����  ��� и����J�      ��  ��� и��I��     �o��G�]z  �E� @�rΓ�7      ��]�vm��  F�� ��	�     �allL� @��  4N�     ���@� @��  � p     耪����  �h� �8�     ���k� h�� ��      �s� �(�;  %�     : ����  F�� ��UU%p     � � h�� ��      �R� �(�;  ��9�     �A� @��  � p     ���  0Z�  � p     �� h�� ��      �R� �(�;  %�     : 缿�  F�� ����      ��;  M� и���      �s� �(�;  �s�     �3��  �h� P��     ��'J�  `t� (A�     ����S�7  0:�  � p     �]�v	� h�� ��U1^z      [3���  ��� ШÇTz      [SU��  4F� @�RJ��7      �u9g�;  �� �(�;     @������  ��� Ш��1�;     @��� @��  4*�,p     萔�� ��� h��     �C\p �Iw  �;     @�� h�� ���)=      ��K)�/� ��!p �i�      pO��^  #p �Q)���      �'w  #p �iw     �n� ��;  ���Z�     �-w  #p �Q)%�;     @����  4F� @��      �s� ��;  M�     t�� ��� hTJI�     �-{""� �h� Ш���      �R-..�;  !p �Q)���      �7u]O��  �h� �4�=      :&�,p �w  �&p     ��;  M� �4�;     @�� h�� �F���      ������  �h� Ш���     �{\p �w  �6Qz       �&�,p �w  ��;     @�� h�� ��	�     �G� @#�  4M�     �=w  !p �iw     ���9� h�� �&��      �"p �w  3333Qz      ���*�;  �� И~�?^z      �.�,p �w  SU��     ���  4B� @c�      �%p �w  �$p     �&�;  �� И��M�;     @7	� h�� �Ƥ�&Jo      `[�  4B� @cRJ.�     t�� �F� h��     ����  �h� И����      ؖ=�  0�  4��k�;     @7�N�>=Vz  >�;  �I)�*�     ��y�W�Ko  ��'p �1w     �����w  �N� @cr�~l%     @GUU%p `��  4�w     ��J)M��  ��O� @c��     tTJ�w  �N� @c\p     �4�;  C'p �19��      ؞�` p `��  4�w     ��J)	� :�;  �I)��     �]w  �N� @cr�.�     t��  4A� @��      �%p `��  4�w     ���Z� ��	� hLJI�     �Q)%�;  C'p �1)���      �6�;  C'p �19g�     �K� ��	� h��     ��RJ�Ko  ��'p �Iw  ��ha    IDAT   �����w  �N� @��      �R�(� ��� ����Jo      `�\p `��  4&��;     @w	� :�;  M�     t�� ��� �$�;     @G���  �� �&	�     :*�,p `��  4i��       �M� ��	� h��      �%p `��  4I�     �]w  �N� @��      �%p `��  4i��       �M� ��	� hJ?|�	     �ew  ��_z��Z^^���z����ґ�����@UU�1Q����R*��-�@D��Ǜ)�A�y="�kq3���s^����N (f}}�������g      �MUUM-//���; �aUJi<�<����kWD�RJ�rν��w5"���=�9窪V#�f]�k?��r���^�wq0\��_��K�w�"��}�K_ZJ)=]����HD����"b|0DDD�9""RJ?�1�u���V?       �v9�^���Z 5��~x�c�1��v����v㻼���"���nD�\U՟���W~�W�7�yT�w�o��o���깈x6">�r��  �w�      �)�9g��Q2O�������:""���W#�ň��񍺮������_����6����Ω�ҧ"��\D�� �j���     ���ATUUz @������^UU,//�DğD���9��~��^,����[�{��{677&��3񩈘+�	 �K�d     ��s� �f#��"��RJ���|!"��s�r����������:A�~��[�����?�s��`0�k)��қ  ��v     t�`0(= �K�"�SJ�86�����R�������7~�7^/=�������9��9����l���G  ;@�     �}�� `��"�r�?���������?�9��]�v��_��_�Rz\���#"眖��2��Ku]����(�	 �A�s����}�eg]�߳ϝ	I�$Pe����ش�VQ���"(-��ը���ҁ{�3#Jr@��9�d���j��"�6`*��,|c�l�4�,�$& M($s3q^�~�G��I2/����}���]k��������^��]:      [d�; �XT9��F�s�9r�`0�����f�d3�������������L)}M�<  ��4     ���� 0vgG�����8~�����ѣ���׼����2��<��녈�ќ�9��  ��     ��w ���g)���:�+���[��:����ҡ�6S����_\U՞�h�҈�� 0K�     �Ϟ ���~�h4z�`0xw]�����sK�\M���{����)�+"��J� �E�y      ��= �Fu"�������`����~fqq��5iS]pEľ�����
�       �V��t �Y�����}0�^J銥����4)SYp_�Rzm������\  �0��      �g� ��/�9�`0��N��waa�s�C��T�{������WD��s��� �?��	     �~�Ѩt  "���l4����:�������C�KU:�������*"���v �m&�\:      [d� ��rnJ�ʺ�?9_T:̸�~����r4��/+� �S��	     �~&� lKO�9�w0�nJ駖����t��h���s���F���v �mN�     ����  lk/�9|8�"�J�٬V��������9�_���K� ��rΥ#      �E&� l{��i8~`8>�t��h]�}8^RUխ���Y  X?�<      �Ϟ @k<?����`𓥃l�\� 뵲�����9����Y  �8�     ��w �V9?"���F?�w�ރ��G+&���:��M�� �R�y      ��= �VzY�ӹy����*d=�}�}m,��qQ�,  l��N     ���� �Z�����u�����N�����ڵ�@�����  �u9��      آ�hT:  �����~0����՟��zGJ:�m9���o|����@� `z��     �~�|  ��ڵ돮��'�r2ۮ������s�Λ#�y��  0>&�     ��	�  �!���cǎ}���?�t�G�V�~���)�E�SJg `�L�      h?{>  S�))�?ۿ�w�r�mSp����>����8�t  ��w     ��3� `��WU��~����A���~��;���xL�,  L�i      �g� `*�L)�z���]:H�6(��=)�k�C  &�b'     @��� �ZUJ���`pE� %/����F�J�  4#�\:      [4�JG  `�^7�*�X�}0�.�T�? ���     �~�|  �_�y�`0(6ļH�����"���z  �c�;     @��� 03��u��x����2�te�� �,�<      ��P# �ّR�r0,5}�F��ಔҵM^ ���b'     @�;v�t  ��?��+�����6yM  �w     ���� 0sRD��.x#)��߿���;#����  �~,v     ��= ��ԩ��7����k�b/����\PU�{"b~�� `���	     �~u]��  @9�s������I_k�����]�N���I^        �<C�  f�W��ͽweee�$/2��{�9u:�_��gL�  ���N        h�g��ͽ#�&u��������dR� �]�     گ���  (,����p�<��O������-��I�        (C� �5o�9���ྲ�rAD�fD̍��  ��	�      �g� �5U��k���x�'��zU��y{J���</  �g�     ����  p\J��UU���덵�>֓���w#���<'        �=�u]:  �HJ�[�=�ܥq�sl��`����q� ��b�     @��� ��RJoX뒏�X
��]w�Y����9�� 0},v       �T�����3�����~�ȑ+"�_��\        ��T�u�  lO_}����8N���p8|fD,�!  S�w     ��Sp �TRJ{����z�-ܯ���9�GĎ� `�)�       �T���_�����-�R�}uu�?F�3�r        �Lp ��y���Wn��.�_s�5O�9_��� 0;Lp     h?w  ��u+++l��M܏;֏��7{<  �E�     ����  ����z�f�T�}���ύ���E          �N)���:����{UU�#"m�X        ���. �vHUU]�s�p�|���`��ƍ �l��	     �~�|  ؀��n�m��~�7t"��7z           fKJ�M�^on#�l��~�w�<".�P*  ���s�      l�	�  l�����d#���6�}�F @��;     �4Pp `~f#S��]p��;~0"���H  �<w     ���� �&<u׮]�a�_^W�}mz��l:  3/�T:      [�� �f�_��I?�u�o����o)  3��*     �O� �Mz�Z'���UpO)-n-        0�� ؤ��|���p�����-� `�Y�     ��}  ،�ҿ���g쥟���s�=�H  �2�      ���  �UU���-����\/["  f��N     ��P�u�  �T������)���>77���1�T        @k)� �;:�Ώ���,��S���          ��X�9���S�8���D        Z�w  �����N��)�u]�|2y           �a�쪟�����/�X           f�K����O��I�v�zaD�h$        �urΥ#  �~�u]��d����s�d�y           �a'�?�����Ή�N<           3)��=�~��G���������1�H*           fN������G����{J�I        �Nιt  �DUU/x�{�|#���<  lUJ�t        `�9� ���b��
����9���          �z�`0���xX�����l           f�N|Q=��om.           �,��-'�~��~�7tRJ��|$  fAJ�t        `�y�7��9�⡂�w��8�H$           f�y��v�3���N����          `���겟Xp��Y           �a)������g� ��H)��      ��KG  `�\|�UD�u�]w^D��bq           �UO�ꪫΏX+�>|��0R          ����;w>+b���*          �6��6b���R��e�  0�R��      �i�s. ����k�����f `�)�        ��Rzz�?LpWp          ���+++�"�+
� `�yT%        p_y�uםW���=�t        �6 `R>�UU]�O* ��R*        �ƪ�zR�Rzb�         @;�� ���u��*"�          (�UD\P:           �-���*"�Q�   L��R�        �6�s~\�+        h��s�  L����;           ��㪈xl�           ̼�V9�sK�  `���JG      `��  0A�V)��S  0�,t        g��J)�,� ���        ���*�l�;        �. 0A;���+� ��g�     `:�� `�vTq�t
  �_UU�#      0
�  L��*�t�t
  ���N     ��`� �	:Z圏�N ����	        ���*�l�;  ��     0��  0AG���j�  L?�      ӡ���  �^�W��)  �~
�      ���  ��R�b_, ��g�     `:�� `Rr�_4� �FX�        N'���*"�_�   L?w     ��`� �II)}���ϖ ����	     0��  0)9绪���t  ���N     ��`� �	��J)�Y:  ��B'     �t�� �����4� �FX�        N'�|Wu����J `�)�     L�>  L�h4��ڷo߽�w��  0�,t     �_Jɾ  ��}���[���T�(  L=�      �g� �I�9*"���H)�U�8  L;��        ���W9�O�� ������_     `[3� �	�ˈ�����Y  �v;     �Ϟ  ��s�h�Z���ѣ�DD.� ��f�     ����  0!ynn�ck�}����.	 ��f�     ����  0!���𥈵���[
� `X�        N����P�=���2Y        �60� �	���?N,��L  fAUUg�      ۚ=  &�.�Cw���w��"�`�8  L=�<      �Ϟ  ������_<Tp��z�RJ.�	 �ig�     ����  0�����g����<  ���        �I�ɉ/Vp����� ��Pp     h?{>  �[J��'�~X�}yy�/"�F 0,v     ��=  ��s������7VpO)���F# 0��:�      ��� �����:�9Y����        ���;  �s~�#�{T�}uu��#��F 03:�N�      l��� 0.)�C9�?x�������z��w  ��b'     @�j ���߻������j�k�y  �1
�      �R* �)�R:ig��-�����E��D 0S�     ��w  �!�t����?�g'm�z�C��&�
 ����     �~&� 0u]�{yy���}vʖQJ魓� ��Qp     h?{>  ��)�ꧼ�\\\�����$�  0{L�      h?w  ��o�����Mp�)��O&  ���锎      �)� 0oI)�S}x�;Δ�["���# 0sLp     h?w  ��hUUo=�N{ǹ��xWD�8�H  �$�     �O� �-�����)��3�|���  0�,v     ���F  lEJ���3�����?>�D  ̬�R�      l�=  ��楥�������Ѽf�a  �q�y      ���� ���|i]w�^x��-� `���     �~
�  lҧWWWߵ�/����K/��V��	 �Yf�     ����  �9�_��z����u�q��Ͽ#"n�l(  f��N     ����^  6*�t����������[F�_~�є�U�� ��Sp     h�N�S:  ���^�wd�_�P���O~�/�?��L  �:w     ��3� ������[6r��ZF�^z�(�t��2 ����<     ��P#  6"����/���F���g��}wD|x�� 0��     گ�锎  @{�����=h�R�/"�&� `F)�     ���  �)G�rJiÝ�Mܻ��"�77s,  ��D     �v����� `���~c�s�a����z1"����  �=      �M� �u8�Rڳك7}ǹgϞ��9�a�� 0{Lp     h7w  �$�����Ż6{���8�;�k"��[9  ��w     �vSp �>>??�VN��;��/��hJ�#��V� �l��	     �n�{  8�c�c�_~����[��\ZZ�hJ�ꭞ ����tJG      `<� ��t����Փ��O*w��qeD|b� `zY�     h7�  8�������8�X
�w�>�s�ш��8y  ��O     �v���ԍ  �.Gs�?�����8N6�;���古�^7�� 0}Lp     h7w  N������q�l�w�|SD��8�	 ��0�     ��� x�]x�+�<�X�8{�^=�~8"�0�� 0Lp     h7�=  �����.����8O:�?�ܻw�9�E�X� �~&z      ��'� ��������{�O<������SJWN��  ��O     �v�� ���v���O�������Ɯ�oM��  ��O     �v��^  "�w����4��O�3���:���['u  �ł'     @���͕�  @Y��ܹ�R��&�0ڽ{�}�N�E��I^ �v0�     ����  ̴{�~��ݻ��E&>BsaaᶈxaD�?�k ����     �n�� 0�H)}��={>=�5r���vo����Q� `{��	     �n ̤QD�����MM\���Q�۽1"~,"rS� `{��J     �v�� 0srD��Z�����v�o�9���k �}X�     h7�=  3g_��}s�l�����|]����.  �UU㷟      ����\�  4��nw�-�0Z^^����ĵ (�D     �v�� 0r΃n����.6Bsyyy9"^_��  4ς'     @�yb/ �Lؿ��.��g�۽2缯d  ���     �^UUEJ�t  &(����v���P�O*���WRJ��Kg `��     ��^ �T�)�奥���ˋ�#"���)������  09Y	     �^
�  S�X��'�����Dl��{D���ү��^��� �dX�     h/{=  S��������_)�mSp��XZZ�ú��w�� ��Y�     h�����  �;���n����AN��
�{��e�ΝGćJg `��     ګ��]� �ͻ���|ݞ={n)䑶�]��ݻ�޹s�wD��Jg `|�     ��^ �������maa�s���̶}n��ݻG������)�AD�H\�    IDATU:  [c�     ����m� ��9�s�.//�b� ��-'��hyy���ƈ�t�,  l��V     ��aF  �R�#���۽�т�{DĞ={n9v�س#���Y  �<��      �e� @k�x���g,--�T:�z��A���7"�w8^�s�>"W:  ��     �^ss�� ��"b���t��hݟU.--�+"�6"��t  6F�     ����  �������m+�G�����vo_]]}~D�:"VK� `}<�     ��� Za5"^����M���]:�f���A�^���kWVV���t������ ��yl%     @{)� l{���v�����o�ݻ��q�`0xID\O*	 �S0�     ��� ��;#�U�n���A�ajF�n����է��E���y  x4��      �e� `{I)J)��F�����1�O���E���W_�ku]_?ST� h;��      �e� `����,,,�V:̸MU�����Ż"��~���RJWD�K#"� 0���     ���; ��������vo.dR���~�������K���3s�?��� 0�����     `�)� ����~vqq��K���h---�E<XtND��9�8"� hXUU�R��s�(      l��; @���{"b����M��4e&
�ǭ��}Ɂ�Z���r�?g�� 0K����hT:      �i�  �9����iaaᓥ�4m&�:>�:p������҈xUD\T8 �L���Sp     h!� &��9��r�Yg�e���w�S�L܏[XX�RD������9�����.��F�Y�� L-�      �d�; �D��߫���C�}���ե��3"�~>8p��c�����e���ʦ �.
�      �� 0V7G�;v����Y��~2�:am���Fį��D�Kr�/N)����� �"�      �d� `KF9���RzOD���vo/h�r�yk�8"��`0��ҋr���_V6 @;Y�     h'�<  ��������rο���|O�@m�s����=�x[�׫�9�g���=�������xlр  -��x(     @�ر�t ���K������СC��zu�Pm��	k�h����s��k��꺮����礔.���"�ܢA �!�=      ��> �����9�RU�MUU}�կ~�_��r�`m�s�~?��󶈈^�W���_u�ر����RJO�������'� �L2�     ��<� �AG#�o#�o"�orΟ��O���}��{����Jd�:
��������<⳹��?��ǎ{|J�	)�'�u��qVUU��9?&"Ύ��a
�vw,"��.�9?����D�h���	?D�߯� 3�ȑ#�O*�     ���9�N<8� fI'"��:�:᧳��s�{;"b5">Q #�s(�r�联���u�ň8\U�=9���??77w����{w��;V �LSp/`��sk?  3�.xgD|�      l�[��֟���?�K�  `�U�  0s(      �����P�  L?w  ����      �qw�}�}  &N� �F�-|     �ϑ�8V:  �O� ��=P:       f� �F(� Ш��Lp     h�C�  0� hT�Y�     �eRJ&� �w  �f�     �er��x  h��;  M3�     �eRJ�Jg  `6(� Ш���;     @˘� @S� h��O     ��1� �F(� ШN�c�;     @�b @#� h��W     ��=  �� @�Lp     h�C�  0� h��      �c� �F(� Ш��	�      �c�;  �Pp �Q9g�=      ��  �Pp �Q���w     ��Qp �
�  4j~~^�     �}� h��;  �:��-~     �ϡ�  �
�  4��[o=��9      �C�  h��;  %.      �1� �F(� P�	      -�s�� @#� (�(     @��� �
�  �`     �ERJ��3  0� (���      X?w  ��� @	�J      `������  �lPp ��     Z����7� �F(� P��;     @{�{���  �Pp ��C�      �n�"�. �٠� @	&|      ����  �
�  4.�d�;     @{��  ��Pp ��     �C� ��(� P�	�      �� @c� h\]�&�     �DJ�`�  �w  J0�     �%r�&� �w  J0�     �=� h��;  %��     �K  `v(� и��	�      -�R2� ��(� P��;     @K�u�� @c� (�P�       ��	�  4I� �ƥ�Lp     hw  �� @	&�     �DJ�`�  �w  ��tLp     h���Mp �1
�  4n׮]
�      -�RRp �1
�  4��[o=�J�      ��RJKg  `v(� Pʡ�      8���Lp �1
�  �r�       ���Ç� h��;  ���     �sssKg  `v(� P�	�      �_���~���!  �
�  �b�;  ��ۻ�9ӳ������n�7Yd��,k,Y���@H��D�!eI@BBd�a�r��d�'$�x�v������~� ��C���y��kg�]��޼���.   �w��ҲG  �>�  dq�     �w�  �^�  d�     ��N�   ֋� �,��      �J.� �Tw  ���     й�� �Tw  Rx3     �����  ��;  )�q���     ����;  K%p  ED�     :�Z��� ��"p  ��     ��5� X*�;  )�q�     t."�  ,�� �.�     L���  ��;  )�      �s� �e� �b�ϲ7      �r�5�;  K%p  ��      ������  �z� �b�;     @��qt� ��� ����w     ���� �R	� H�����2f�      ��Ο?�;  K%p  �XJ��=     �:���z�= ��"p  ӝ�      ����  ��;  �>�      �d  `�� ��;     @�"B� ��	� �$p     �Tk�v�  ֏� �Lw     �N��\p `��  d�     t*"\p `��  �i�	�     ��;  K'p  MD�     :w  �N� @�;     @�Zk��7  �~�  ����      <��  d� ��w     �~�� @�;  i�      ���w  �N� @�q�      ��A� ��	� H�;     @����ogo  `�� HSk�     tjcc�w  �N� @�Ǐ�     �Ԯ^��Y�  ֏� �4��̛�      }�[J9� ��� �f{{���Ҳw      �7�  ���  d:*���     �� H!p  ���      |�� �w  �d      ��  �� ��w     ��� H!p  ��     �?w  R� �&p     �� �w  �	�     �#p  �� �T�5�;     @gZkw  R� H�      ��;  )�  �r�     �?�8
� H!p  U�U�     ЙǏ� H!p  ��      �y|�֭;�#  XOw  R��(p     �˭RJ� �z� �j6�	�     �r3{   �K� @���#�;     @_�  �� ��_���     �/w  �� Hu���ǥ���;      �w  �� �+�      �� �F� @�      �� �F� @�      �� �F� @�֚�     �w  �� Hw     �N���  �� ��;     @'�  d� ��w     �~��(p  �� �t����      �֗����do  `}	� H�Zs�     ��.]z�= ��%p  ]�U�     Ё���� ��&p  ]k�V�      Ji����  �z� ��@      ���  �z� ��;     @�  �� ����X�     Ё֚� �Tw  �-�{���;      �]D� H%p ���      ������  �z� Ћ��      ��8�.� �J� @/�      �j�w  R	� ��~�      �u���)p  �� �.��\p     �������#  Xow  z!p     ��z;  ��  t��*p     H�Z� �N� @/�      �"b/{  � �BD�go      Xs.� �N� @/\p     H�Z� �N� @/�      �"B� @:�;  ]��
�     	� �� �.\�z�v)�({     ���q/{  � �E+��&{     ������ @:�;  =��=      `]mnn
� H'p �'w     �/_�|�=  �  �d?{      ��r� �.� ��      	Zkw  � p �'w     �!p �w  z"p     ȱ�=   J� ��;     @�֚�  tA� @O��      ���� ��;  ���)     @�k�  ��;  9::�     $h�ͳ7  @)w  �"p     H0���  tA� @7�ŽR���      k�p�X��  �� �+�      Kۥ���  J� ��;     �r]�   �� ��;     �����  �sw  ��Z�     ,��  tC� @W"B�     �\.� ��;  ]�     ,�� �n� ��8�w     �庖=   >'p �+���     `��� @7�  te�     ��p�X��  �� Е�
�     �g^Ji�#  �sw  �r�ƍ���{�;      �AD̳7  ���  ��z�      �u�Z� ��;  =Zd      Xײ  ���  �h/{      ��p� ��� �Nk�w     ��� ��;  ݉�;     �r\�   O� �#�;     ��� @W�  t��&p     8{����F�  x�� ��D��     ���K)-{  <M� @wj�w     �3��  �,�;  ��q;{     ��k�meo  �g	� ������Rʭ�      +���  �,�;  ��      g("�  tG� @�Zkw     �3�Z���  �%p �Wײ      ��Z��  tG� @�j���      V��|>��  �� Х��<{     �
�*���#  �Yw  z%p     8;�f  ��� Ыk�      V�� �.	� �����     ��� �� �.-�{����;      VQk�r�  x�;  ݊�y�     �UTk�u�  x�;  �j�	�     ����� �.	� �ٵ�      +ho�N�  x�;  =��      ��~�=   ^d�=   ^b�Z+��� /t���rpp�=���ѣ2�c�    �Rk-E� @��  t��6?<<�]������׳g@��Ey��a�    ��/}��R>��  /R�  ���֮eo      X5�V� �� �n	�     N�� �n	� ������Z���      �""������  �"w  z��      �
"��Rv����do �� е����      �
��d�  ��� е��V�     �U�����  �2w  �VkuE     �<��.p �kw  ����     `DD��;  ]� е�l�MV     �S�$p�8{  ��� ��=z��'_�	     �[���������  /#p �k7nܸ�;      V�/J)-{  ��� �)pI     �-DD��^��  �"p �{�֭�      S�����  �*w  ��Z�${     ���ZK)���  �*w  �7�k"      o��Zj�>s �{w  �7�k"      o!"������;  �U�  tocc�W�=     `�"�J)c�  x�;  ݻr��^��a�     ������  pw  ��E�N�     �)�����G�;  �$�  L�V�      �)� 0%w  &�����      Smss�g�;  �$�  L�0���      0E����u;{  ��� ���yDdo      ��Z�G�  ��  L�0��     ���(�0|��  NJ� �$���Ok���w      LI����x1{  ��� ��8��ne�      ��Zk���d�  ��� 0�q�     �)�����ٹ��  NJ� �d��Q�     �)q� ��� 0%��     �$"��Z��  ^�: �ɨ�
�     N���*�w  ��P 0��엵�1{     ��Z˹s�~��  ^�� �����zW�w      LA�u�ʕ+��;  �u� ��a~��     `
�a�Q�  x]w  �惈��      еZk)��w�  x]w  &����'o�     ���w  &G �������     ��axx���w  ��R 0)����Z���      =����ҥK��w  ��� 05���Q�     �^ED��~/{  �	�;  �DD�     �.�P"���;  �M� ����Ok�(     �<�0���d�  �7�
 `���     <_D\��緲w  ��P 09���G�0<��     Л�(����  oJ� ��\�x�q����      ����R���  oJ� �$E�k�8     �ak����  oJ �$��~$p     �]�0|o>�?��  oJ �$���'_�	     @)��g'���  oC� �$]�v�r�u?{     @/�a(�n�  xw  ��E�k�H     PJ)�ֽ���f�  ��� `���     �����RJ��  oC �d�����0d�      H7��J)�;�;  �m	� ������#� {     @�Z��W����w  ��� 0e���Z=�     ��Z�a�ǋ/>��  oK	 ��E�{�0d�      H�䳒�d�  �� p `�Zk��;     ��f���Rʻ�;  �4(�  ����݋�0lg�      �Pk-�͝����[  �4� ��VJ��'_�	     �Vf�Y���g�  ��"p `���     XG�0�r{{��;  �� X��� {     �2=������o� �� p `�vvv�R��V��     ��������7�w  �iR  �*�9�Ͳ7      ,E����wׯ__do ��$p `%Dķ�a���     `f��8���d�  ��&p `%���܏����#.     ��"��f�o���}��  N�� ��Qk��l6˞     p�666Jk�w  �Y� �2���{��̥     `eED���������-  p�  ���Z�+W�    �U���qw�?��  gE� �J�����l6�u�     ����c�  �IDAT6C��/���v�  8+w  V�q��/�a��     p�Ν;�㝝����  gI� ��������s��-{     �i����Mk�OJ)��[  �,	� XE-"�l6���     �f��݈���b�i�  8kw  V����s���iq�     ���l�����{{{?��  � p `e���~kss�K)7��      ��Z��l������������{  `Yf�  �,-�*�|�TJ���X=<x��͛���:�[Jy�=  ���ZJN�Ν���͎�����f��8����儍Gk���x*��g�M�^��~ "�k��[��Q)�=��G���q)�w��a~�5#�?���Xk�=����s�  �v���R�y�L    IEND�B`�PK
     ���Z'�Y��  �  /   images/4bf63cb1-3675-4452-8ab6-1403298522d5.png�PNG

   IHDR   d      X�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  SIDATx���KA�_�&�Ҕj�PZL-1����?�7O=x��[�ދ'�{�xl=x#"�P"�ɖ�T�[b�&���ݢv��xa��o�;o�f&
I ��ё��v��F��5�M������Yj�ۧ�����ZZZ��v�����$��\�v�T�)�Q�Z���?�;r�V�B�x�1E����� &M6���������FM�0��UUu���[�;<<$��K�Z�L���B�@�LF/_7Ft�o}<YB��.��Ȉ�8��p�\�b�hY��|>D�A=�\����l!�>����=�����y�ϐ!v�[V�������ѓ�=��a��ò���;�\��)�mr.�&�277'�A,C�d�����ƉpF��F)�uI�
f�`���(_���X��N�ǐ�v�����4�q$����"�q�	T���.�[�$�F���E��:MdW���a��n��4�'�b�to���f�����<��.�1L� �=�%n ���r�F�I�wQR�V!��{�G"[��Zbh_+���Ol3$����%��;�'���������(Ϥ'�0�j�����U�99��Xf{Ƕk�Cv�8����
�����v� ;;;����W��t)�x�D�ֱLmll ��PX���ښ^����.�P̂(p$mP!��/eqqQh��!Fk�\��jX� 8.1�d�"��{�n��Il�~�&#��r���>�t�z�JE���>��-��ޞ^�n�a<I��+nDE#E������O�[V�0��T*u�pZl�k'���UV�R1�n�y0q�<��>���$���I�"�t}�4���������J�u�    IEND�B`�PK 
     ���Z�ަ���  ��                   cirkitFile.jsonPK 
     ���Z                        ̯  jsons/PK 
     ���Z71��8  �8               �  jsons/user_defined.jsonPK 
     ���Z                        ��  images/PK 
     ���Z�?.�� � /             ��  images/1fa09ac9-b6db-4b4a-b77c-89392a61857d.pngPK 
     ���Z�ȽF �F /             , images/c5aba2f5-4dea-4d75-9bc6-8c6f78bbb1f3.pngPK 
     ���Zv'ON��  ��  /             6H images/0755f9ac-cddf-41fa-8c34-4d71983a54be.pngPK 
     ���Z�����  ��  /             _1 images/2abdabbf-059f-44b6-b68f-d45f0cb3c7dc.pngPK 
     ���Zq���W W /             � images/7c9bed20-c7d7-43dc-b689-820375f46db8.pngPK 
     ���Z$�3  3  /             �q images/7ade412b-fa94-47ea-987a-d6c9baa14438.pngPK 
     ���Z��F�} �} /             r� images/b63deb06-c33f-4ae3-8f73-25229955b1c1.pngPK 
     ���Z���  �  /             � images/a5640015-ff5c-4848-bb8b-6d4b42e5489b.pngPK 
     ���Z	��} } /             � images/bbfae99c-8036-4c5e-89fd-a87441410720.pngPK 
     ���Zd��   �   /             @� images/a262aa33-74c4-460b-b0ad-c746896f6744.pngPK 
     ���Z"1^FHo Ho /             � images/4efcf596-32b1-4e3b-9735-2bd5fa764fde.pngPK 
     ���Z��n  n  /             �' images/a46afb92-29a7-4c70-92b4-1e1235f7410a.pngPK 
     ���Z�&�y`  y`  /             h@ images/8c2f1315-cf23-4ba8-a920-becb97f13280.pngPK 
     ���Z�����  �  /             .� images/6fc4b800-efc3-4a5d-827d-9566cfd108b3.pngPK 
     ���Z
�8b  8b  /             h� images/a7e3301e-fb46-458d-916f-a05c0bde95f4.pngPK 
     ���Z'�Y��  �  /             � images/4bf63cb1-3675-4452-8ab6-1403298522d5.pngPK      �      